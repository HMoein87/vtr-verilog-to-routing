

/*
 *
 * RAW Benchmark Suite main defines
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz 

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/jacobi/src/library.v,v 1.5 1997/08/09 05:57:41 jbabb Exp $
 *
 * Library for Jacobi benchmark
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 * This is the behavioral verilog library for this benchmark.
 * By convention, all module names start with the benchmark name.
 * All top-level modules must have the global connections:
 *   Clk, Reset, RD, WR, Addr, DataIn, DataOut
 * Modules may also have any number of local connections or
 * sub-modules without restriction.
 *
 */


/* The basic array node */

module Jacobi_Node (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		    ScanIn, ScanOut, ScanEnable,
		    Id, Enable, NorthIn, SouthIn, EastIn, WestIn, Out);
   
   parameter WIDTH    = 8,
	     IDWIDTH  = 8,
	     BOUNDARY = 0,
	     SCAN     = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;   


   /* local connections */
   
   input			 Enable;
   input [IDWIDTH-1:0]		 Id;
   input [WIDTH-1:0]		 NorthIn,SouthIn,EastIn,WestIn;
   output [WIDTH-1:0]		 Out;
   
   reg [WIDTH-1:0]		 Out;
   
   
   /* support reading of the node data value (non-scan only) */
   
   assign DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out: `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;

   
   always @(posedge Clk)
      begin	

	 
	 /* reset will initialize the entire array to zero */
	 
	 if (Reset)
	    Out=0;	 


	 /* support scan in */

	 else if (SCAN && ScanEnable)
	    Out=ScanIn[WIDTH-1:0];
	 

	 /* support writing of the node data value (non-scan only) */
	 
	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0]==Id))
	    Out=DataIn[WIDTH-1:0];
	 

	 /* for non-boundary nodes, do the Jacobi computation when enabled */
	 
	 else if (!BOUNDARY && Enable)
	    Out=(NorthIn+SouthIn+EastIn+WestIn) >> 2;

      end
endmodule


/* 
 * A control module to count iterations.
 *
 * Writing to Address==ID will set a counter.
 *
 * The other Jacobi nodes will be enabled by this module when 
 * count is greater than zero.
 *
 * The counter will decrement every cycle down to zero.
 *
 * This module also handles scan control.
 */

module Jacobi_Control (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		       ScanIn, ScanOut, ScanEnable,
		       Id,ScanId,Enable);
   
   parameter WIDTH   = 8,
	     CWIDTH  = 8,
	     IDWIDTH = 8,
	     SCAN    = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [IDWIDTH-1:0]		 ScanId;
   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;   


   /* local connections */
   
   input [IDWIDTH-1:0]		 Id;
   output			 Enable;
   
   
   /* a register for the counter and scan */

   reg [CWIDTH-1:0]		 count;
   reg [WIDTH-1:0]		 ScanReg;

   
   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? count:
      (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;
   
   
   /* enable when count is active */
   
   assign Enable = !(count==0);

   
   always @(posedge Clk)
      begin

	 
	 /* store current scan output */

	 ScanReg=ScanIn;


	 /* Logic to reset, write, and decrement the counter */
	 
	 if (Reset)
	    count=0;
	 else if (WR && (Addr[IDWIDTH-1:0]==Id))
	    count=DataIn[CWIDTH-1:0];
	 else if(count) 
	    count=count-1;
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [7:0] nOut0_0;
wire [7:0] nScanOut0;
wire [7:0] nOut0_1;
wire [7:0] nScanOut1;
wire [7:0] nOut0_2;
wire [7:0] nScanOut2;
wire [7:0] nOut0_3;
wire [7:0] nScanOut3;
wire [7:0] nOut0_4;
wire [7:0] nScanOut4;
wire [7:0] nOut0_5;
wire [7:0] nScanOut5;
wire [7:0] nOut0_6;
wire [7:0] nScanOut6;
wire [7:0] nOut0_7;
wire [7:0] nScanOut7;
wire [7:0] nOut0_8;
wire [7:0] nScanOut8;
wire [7:0] nOut0_9;
wire [7:0] nScanOut9;
wire [7:0] nOut0_10;
wire [7:0] nScanOut10;
wire [7:0] nOut0_11;
wire [7:0] nScanOut11;
wire [7:0] nOut0_12;
wire [7:0] nScanOut12;
wire [7:0] nOut0_13;
wire [7:0] nScanOut13;
wire [7:0] nOut0_14;
wire [7:0] nScanOut14;
wire [7:0] nOut0_15;
wire [7:0] nScanOut15;
wire [7:0] nOut0_16;
wire [7:0] nScanOut16;
wire [7:0] nOut0_17;
wire [7:0] nScanOut17;
wire [7:0] nOut0_18;
wire [7:0] nScanOut18;
wire [7:0] nOut0_19;
wire [7:0] nScanOut19;
wire [7:0] nOut0_20;
wire [7:0] nScanOut20;
wire [7:0] nOut0_21;
wire [7:0] nScanOut21;
wire [7:0] nOut0_22;
wire [7:0] nScanOut22;
wire [7:0] nOut0_23;
wire [7:0] nScanOut23;
wire [7:0] nOut0_24;
wire [7:0] nScanOut24;
wire [7:0] nOut0_25;
wire [7:0] nScanOut25;
wire [7:0] nOut0_26;
wire [7:0] nScanOut26;
wire [7:0] nOut0_27;
wire [7:0] nScanOut27;
wire [7:0] nOut0_28;
wire [7:0] nScanOut28;
wire [7:0] nOut0_29;
wire [7:0] nScanOut29;
wire [7:0] nOut0_30;
wire [7:0] nScanOut30;
wire [7:0] nOut0_31;
wire [7:0] nScanOut31;
wire [7:0] nOut0_32;
wire [7:0] nScanOut32;
wire [7:0] nOut0_33;
wire [7:0] nScanOut33;
wire [7:0] nOut0_34;
wire [7:0] nScanOut34;
wire [7:0] nOut0_35;
wire [7:0] nScanOut35;
wire [7:0] nOut0_36;
wire [7:0] nScanOut36;
wire [7:0] nOut0_37;
wire [7:0] nScanOut37;
wire [7:0] nOut0_38;
wire [7:0] nScanOut38;
wire [7:0] nOut0_39;
wire [7:0] nScanOut39;
wire [7:0] nOut0_40;
wire [7:0] nScanOut40;
wire [7:0] nOut0_41;
wire [7:0] nScanOut41;
wire [7:0] nOut0_42;
wire [7:0] nScanOut42;
wire [7:0] nOut0_43;
wire [7:0] nScanOut43;
wire [7:0] nOut0_44;
wire [7:0] nScanOut44;
wire [7:0] nOut0_45;
wire [7:0] nScanOut45;
wire [7:0] nOut0_46;
wire [7:0] nScanOut46;
wire [7:0] nOut0_47;
wire [7:0] nScanOut47;
wire [7:0] nOut0_48;
wire [7:0] nScanOut48;
wire [7:0] nOut0_49;
wire [7:0] nScanOut49;
wire [7:0] nOut0_50;
wire [7:0] nScanOut50;
wire [7:0] nOut0_51;
wire [7:0] nScanOut51;
wire [7:0] nOut0_52;
wire [7:0] nScanOut52;
wire [7:0] nOut0_53;
wire [7:0] nScanOut53;
wire [7:0] nOut0_54;
wire [7:0] nScanOut54;
wire [7:0] nOut0_55;
wire [7:0] nScanOut55;
wire [7:0] nOut0_56;
wire [7:0] nScanOut56;
wire [7:0] nOut0_57;
wire [7:0] nScanOut57;
wire [7:0] nOut0_58;
wire [7:0] nScanOut58;
wire [7:0] nOut0_59;
wire [7:0] nScanOut59;
wire [7:0] nOut0_60;
wire [7:0] nScanOut60;
wire [7:0] nOut0_61;
wire [7:0] nScanOut61;
wire [7:0] nOut0_62;
wire [7:0] nScanOut62;
wire [7:0] nOut0_63;
wire [7:0] nScanOut63;
wire [7:0] nOut1_0;
wire [7:0] nScanOut64;
wire [7:0] nOut1_1;
wire [7:0] nScanOut65;
wire [7:0] nOut1_2;
wire [7:0] nScanOut66;
wire [7:0] nOut1_3;
wire [7:0] nScanOut67;
wire [7:0] nOut1_4;
wire [7:0] nScanOut68;
wire [7:0] nOut1_5;
wire [7:0] nScanOut69;
wire [7:0] nOut1_6;
wire [7:0] nScanOut70;
wire [7:0] nOut1_7;
wire [7:0] nScanOut71;
wire [7:0] nOut1_8;
wire [7:0] nScanOut72;
wire [7:0] nOut1_9;
wire [7:0] nScanOut73;
wire [7:0] nOut1_10;
wire [7:0] nScanOut74;
wire [7:0] nOut1_11;
wire [7:0] nScanOut75;
wire [7:0] nOut1_12;
wire [7:0] nScanOut76;
wire [7:0] nOut1_13;
wire [7:0] nScanOut77;
wire [7:0] nOut1_14;
wire [7:0] nScanOut78;
wire [7:0] nOut1_15;
wire [7:0] nScanOut79;
wire [7:0] nOut1_16;
wire [7:0] nScanOut80;
wire [7:0] nOut1_17;
wire [7:0] nScanOut81;
wire [7:0] nOut1_18;
wire [7:0] nScanOut82;
wire [7:0] nOut1_19;
wire [7:0] nScanOut83;
wire [7:0] nOut1_20;
wire [7:0] nScanOut84;
wire [7:0] nOut1_21;
wire [7:0] nScanOut85;
wire [7:0] nOut1_22;
wire [7:0] nScanOut86;
wire [7:0] nOut1_23;
wire [7:0] nScanOut87;
wire [7:0] nOut1_24;
wire [7:0] nScanOut88;
wire [7:0] nOut1_25;
wire [7:0] nScanOut89;
wire [7:0] nOut1_26;
wire [7:0] nScanOut90;
wire [7:0] nOut1_27;
wire [7:0] nScanOut91;
wire [7:0] nOut1_28;
wire [7:0] nScanOut92;
wire [7:0] nOut1_29;
wire [7:0] nScanOut93;
wire [7:0] nOut1_30;
wire [7:0] nScanOut94;
wire [7:0] nOut1_31;
wire [7:0] nScanOut95;
wire [7:0] nOut1_32;
wire [7:0] nScanOut96;
wire [7:0] nOut1_33;
wire [7:0] nScanOut97;
wire [7:0] nOut1_34;
wire [7:0] nScanOut98;
wire [7:0] nOut1_35;
wire [7:0] nScanOut99;
wire [7:0] nOut1_36;
wire [7:0] nScanOut100;
wire [7:0] nOut1_37;
wire [7:0] nScanOut101;
wire [7:0] nOut1_38;
wire [7:0] nScanOut102;
wire [7:0] nOut1_39;
wire [7:0] nScanOut103;
wire [7:0] nOut1_40;
wire [7:0] nScanOut104;
wire [7:0] nOut1_41;
wire [7:0] nScanOut105;
wire [7:0] nOut1_42;
wire [7:0] nScanOut106;
wire [7:0] nOut1_43;
wire [7:0] nScanOut107;
wire [7:0] nOut1_44;
wire [7:0] nScanOut108;
wire [7:0] nOut1_45;
wire [7:0] nScanOut109;
wire [7:0] nOut1_46;
wire [7:0] nScanOut110;
wire [7:0] nOut1_47;
wire [7:0] nScanOut111;
wire [7:0] nOut1_48;
wire [7:0] nScanOut112;
wire [7:0] nOut1_49;
wire [7:0] nScanOut113;
wire [7:0] nOut1_50;
wire [7:0] nScanOut114;
wire [7:0] nOut1_51;
wire [7:0] nScanOut115;
wire [7:0] nOut1_52;
wire [7:0] nScanOut116;
wire [7:0] nOut1_53;
wire [7:0] nScanOut117;
wire [7:0] nOut1_54;
wire [7:0] nScanOut118;
wire [7:0] nOut1_55;
wire [7:0] nScanOut119;
wire [7:0] nOut1_56;
wire [7:0] nScanOut120;
wire [7:0] nOut1_57;
wire [7:0] nScanOut121;
wire [7:0] nOut1_58;
wire [7:0] nScanOut122;
wire [7:0] nOut1_59;
wire [7:0] nScanOut123;
wire [7:0] nOut1_60;
wire [7:0] nScanOut124;
wire [7:0] nOut1_61;
wire [7:0] nScanOut125;
wire [7:0] nOut1_62;
wire [7:0] nScanOut126;
wire [7:0] nOut1_63;
wire [7:0] nScanOut127;
wire [7:0] nOut2_0;
wire [7:0] nScanOut128;
wire [7:0] nOut2_1;
wire [7:0] nScanOut129;
wire [7:0] nOut2_2;
wire [7:0] nScanOut130;
wire [7:0] nOut2_3;
wire [7:0] nScanOut131;
wire [7:0] nOut2_4;
wire [7:0] nScanOut132;
wire [7:0] nOut2_5;
wire [7:0] nScanOut133;
wire [7:0] nOut2_6;
wire [7:0] nScanOut134;
wire [7:0] nOut2_7;
wire [7:0] nScanOut135;
wire [7:0] nOut2_8;
wire [7:0] nScanOut136;
wire [7:0] nOut2_9;
wire [7:0] nScanOut137;
wire [7:0] nOut2_10;
wire [7:0] nScanOut138;
wire [7:0] nOut2_11;
wire [7:0] nScanOut139;
wire [7:0] nOut2_12;
wire [7:0] nScanOut140;
wire [7:0] nOut2_13;
wire [7:0] nScanOut141;
wire [7:0] nOut2_14;
wire [7:0] nScanOut142;
wire [7:0] nOut2_15;
wire [7:0] nScanOut143;
wire [7:0] nOut2_16;
wire [7:0] nScanOut144;
wire [7:0] nOut2_17;
wire [7:0] nScanOut145;
wire [7:0] nOut2_18;
wire [7:0] nScanOut146;
wire [7:0] nOut2_19;
wire [7:0] nScanOut147;
wire [7:0] nOut2_20;
wire [7:0] nScanOut148;
wire [7:0] nOut2_21;
wire [7:0] nScanOut149;
wire [7:0] nOut2_22;
wire [7:0] nScanOut150;
wire [7:0] nOut2_23;
wire [7:0] nScanOut151;
wire [7:0] nOut2_24;
wire [7:0] nScanOut152;
wire [7:0] nOut2_25;
wire [7:0] nScanOut153;
wire [7:0] nOut2_26;
wire [7:0] nScanOut154;
wire [7:0] nOut2_27;
wire [7:0] nScanOut155;
wire [7:0] nOut2_28;
wire [7:0] nScanOut156;
wire [7:0] nOut2_29;
wire [7:0] nScanOut157;
wire [7:0] nOut2_30;
wire [7:0] nScanOut158;
wire [7:0] nOut2_31;
wire [7:0] nScanOut159;
wire [7:0] nOut2_32;
wire [7:0] nScanOut160;
wire [7:0] nOut2_33;
wire [7:0] nScanOut161;
wire [7:0] nOut2_34;
wire [7:0] nScanOut162;
wire [7:0] nOut2_35;
wire [7:0] nScanOut163;
wire [7:0] nOut2_36;
wire [7:0] nScanOut164;
wire [7:0] nOut2_37;
wire [7:0] nScanOut165;
wire [7:0] nOut2_38;
wire [7:0] nScanOut166;
wire [7:0] nOut2_39;
wire [7:0] nScanOut167;
wire [7:0] nOut2_40;
wire [7:0] nScanOut168;
wire [7:0] nOut2_41;
wire [7:0] nScanOut169;
wire [7:0] nOut2_42;
wire [7:0] nScanOut170;
wire [7:0] nOut2_43;
wire [7:0] nScanOut171;
wire [7:0] nOut2_44;
wire [7:0] nScanOut172;
wire [7:0] nOut2_45;
wire [7:0] nScanOut173;
wire [7:0] nOut2_46;
wire [7:0] nScanOut174;
wire [7:0] nOut2_47;
wire [7:0] nScanOut175;
wire [7:0] nOut2_48;
wire [7:0] nScanOut176;
wire [7:0] nOut2_49;
wire [7:0] nScanOut177;
wire [7:0] nOut2_50;
wire [7:0] nScanOut178;
wire [7:0] nOut2_51;
wire [7:0] nScanOut179;
wire [7:0] nOut2_52;
wire [7:0] nScanOut180;
wire [7:0] nOut2_53;
wire [7:0] nScanOut181;
wire [7:0] nOut2_54;
wire [7:0] nScanOut182;
wire [7:0] nOut2_55;
wire [7:0] nScanOut183;
wire [7:0] nOut2_56;
wire [7:0] nScanOut184;
wire [7:0] nOut2_57;
wire [7:0] nScanOut185;
wire [7:0] nOut2_58;
wire [7:0] nScanOut186;
wire [7:0] nOut2_59;
wire [7:0] nScanOut187;
wire [7:0] nOut2_60;
wire [7:0] nScanOut188;
wire [7:0] nOut2_61;
wire [7:0] nScanOut189;
wire [7:0] nOut2_62;
wire [7:0] nScanOut190;
wire [7:0] nOut2_63;
wire [7:0] nScanOut191;
wire [7:0] nOut3_0;
wire [7:0] nScanOut192;
wire [7:0] nOut3_1;
wire [7:0] nScanOut193;
wire [7:0] nOut3_2;
wire [7:0] nScanOut194;
wire [7:0] nOut3_3;
wire [7:0] nScanOut195;
wire [7:0] nOut3_4;
wire [7:0] nScanOut196;
wire [7:0] nOut3_5;
wire [7:0] nScanOut197;
wire [7:0] nOut3_6;
wire [7:0] nScanOut198;
wire [7:0] nOut3_7;
wire [7:0] nScanOut199;
wire [7:0] nOut3_8;
wire [7:0] nScanOut200;
wire [7:0] nOut3_9;
wire [7:0] nScanOut201;
wire [7:0] nOut3_10;
wire [7:0] nScanOut202;
wire [7:0] nOut3_11;
wire [7:0] nScanOut203;
wire [7:0] nOut3_12;
wire [7:0] nScanOut204;
wire [7:0] nOut3_13;
wire [7:0] nScanOut205;
wire [7:0] nOut3_14;
wire [7:0] nScanOut206;
wire [7:0] nOut3_15;
wire [7:0] nScanOut207;
wire [7:0] nOut3_16;
wire [7:0] nScanOut208;
wire [7:0] nOut3_17;
wire [7:0] nScanOut209;
wire [7:0] nOut3_18;
wire [7:0] nScanOut210;
wire [7:0] nOut3_19;
wire [7:0] nScanOut211;
wire [7:0] nOut3_20;
wire [7:0] nScanOut212;
wire [7:0] nOut3_21;
wire [7:0] nScanOut213;
wire [7:0] nOut3_22;
wire [7:0] nScanOut214;
wire [7:0] nOut3_23;
wire [7:0] nScanOut215;
wire [7:0] nOut3_24;
wire [7:0] nScanOut216;
wire [7:0] nOut3_25;
wire [7:0] nScanOut217;
wire [7:0] nOut3_26;
wire [7:0] nScanOut218;
wire [7:0] nOut3_27;
wire [7:0] nScanOut219;
wire [7:0] nOut3_28;
wire [7:0] nScanOut220;
wire [7:0] nOut3_29;
wire [7:0] nScanOut221;
wire [7:0] nOut3_30;
wire [7:0] nScanOut222;
wire [7:0] nOut3_31;
wire [7:0] nScanOut223;
wire [7:0] nOut3_32;
wire [7:0] nScanOut224;
wire [7:0] nOut3_33;
wire [7:0] nScanOut225;
wire [7:0] nOut3_34;
wire [7:0] nScanOut226;
wire [7:0] nOut3_35;
wire [7:0] nScanOut227;
wire [7:0] nOut3_36;
wire [7:0] nScanOut228;
wire [7:0] nOut3_37;
wire [7:0] nScanOut229;
wire [7:0] nOut3_38;
wire [7:0] nScanOut230;
wire [7:0] nOut3_39;
wire [7:0] nScanOut231;
wire [7:0] nOut3_40;
wire [7:0] nScanOut232;
wire [7:0] nOut3_41;
wire [7:0] nScanOut233;
wire [7:0] nOut3_42;
wire [7:0] nScanOut234;
wire [7:0] nOut3_43;
wire [7:0] nScanOut235;
wire [7:0] nOut3_44;
wire [7:0] nScanOut236;
wire [7:0] nOut3_45;
wire [7:0] nScanOut237;
wire [7:0] nOut3_46;
wire [7:0] nScanOut238;
wire [7:0] nOut3_47;
wire [7:0] nScanOut239;
wire [7:0] nOut3_48;
wire [7:0] nScanOut240;
wire [7:0] nOut3_49;
wire [7:0] nScanOut241;
wire [7:0] nOut3_50;
wire [7:0] nScanOut242;
wire [7:0] nOut3_51;
wire [7:0] nScanOut243;
wire [7:0] nOut3_52;
wire [7:0] nScanOut244;
wire [7:0] nOut3_53;
wire [7:0] nScanOut245;
wire [7:0] nOut3_54;
wire [7:0] nScanOut246;
wire [7:0] nOut3_55;
wire [7:0] nScanOut247;
wire [7:0] nOut3_56;
wire [7:0] nScanOut248;
wire [7:0] nOut3_57;
wire [7:0] nScanOut249;
wire [7:0] nOut3_58;
wire [7:0] nScanOut250;
wire [7:0] nOut3_59;
wire [7:0] nScanOut251;
wire [7:0] nOut3_60;
wire [7:0] nScanOut252;
wire [7:0] nOut3_61;
wire [7:0] nScanOut253;
wire [7:0] nOut3_62;
wire [7:0] nScanOut254;
wire [7:0] nOut3_63;
wire [7:0] nScanOut255;
wire [7:0] nOut4_0;
wire [7:0] nScanOut256;
wire [7:0] nOut4_1;
wire [7:0] nScanOut257;
wire [7:0] nOut4_2;
wire [7:0] nScanOut258;
wire [7:0] nOut4_3;
wire [7:0] nScanOut259;
wire [7:0] nOut4_4;
wire [7:0] nScanOut260;
wire [7:0] nOut4_5;
wire [7:0] nScanOut261;
wire [7:0] nOut4_6;
wire [7:0] nScanOut262;
wire [7:0] nOut4_7;
wire [7:0] nScanOut263;
wire [7:0] nOut4_8;
wire [7:0] nScanOut264;
wire [7:0] nOut4_9;
wire [7:0] nScanOut265;
wire [7:0] nOut4_10;
wire [7:0] nScanOut266;
wire [7:0] nOut4_11;
wire [7:0] nScanOut267;
wire [7:0] nOut4_12;
wire [7:0] nScanOut268;
wire [7:0] nOut4_13;
wire [7:0] nScanOut269;
wire [7:0] nOut4_14;
wire [7:0] nScanOut270;
wire [7:0] nOut4_15;
wire [7:0] nScanOut271;
wire [7:0] nOut4_16;
wire [7:0] nScanOut272;
wire [7:0] nOut4_17;
wire [7:0] nScanOut273;
wire [7:0] nOut4_18;
wire [7:0] nScanOut274;
wire [7:0] nOut4_19;
wire [7:0] nScanOut275;
wire [7:0] nOut4_20;
wire [7:0] nScanOut276;
wire [7:0] nOut4_21;
wire [7:0] nScanOut277;
wire [7:0] nOut4_22;
wire [7:0] nScanOut278;
wire [7:0] nOut4_23;
wire [7:0] nScanOut279;
wire [7:0] nOut4_24;
wire [7:0] nScanOut280;
wire [7:0] nOut4_25;
wire [7:0] nScanOut281;
wire [7:0] nOut4_26;
wire [7:0] nScanOut282;
wire [7:0] nOut4_27;
wire [7:0] nScanOut283;
wire [7:0] nOut4_28;
wire [7:0] nScanOut284;
wire [7:0] nOut4_29;
wire [7:0] nScanOut285;
wire [7:0] nOut4_30;
wire [7:0] nScanOut286;
wire [7:0] nOut4_31;
wire [7:0] nScanOut287;
wire [7:0] nOut4_32;
wire [7:0] nScanOut288;
wire [7:0] nOut4_33;
wire [7:0] nScanOut289;
wire [7:0] nOut4_34;
wire [7:0] nScanOut290;
wire [7:0] nOut4_35;
wire [7:0] nScanOut291;
wire [7:0] nOut4_36;
wire [7:0] nScanOut292;
wire [7:0] nOut4_37;
wire [7:0] nScanOut293;
wire [7:0] nOut4_38;
wire [7:0] nScanOut294;
wire [7:0] nOut4_39;
wire [7:0] nScanOut295;
wire [7:0] nOut4_40;
wire [7:0] nScanOut296;
wire [7:0] nOut4_41;
wire [7:0] nScanOut297;
wire [7:0] nOut4_42;
wire [7:0] nScanOut298;
wire [7:0] nOut4_43;
wire [7:0] nScanOut299;
wire [7:0] nOut4_44;
wire [7:0] nScanOut300;
wire [7:0] nOut4_45;
wire [7:0] nScanOut301;
wire [7:0] nOut4_46;
wire [7:0] nScanOut302;
wire [7:0] nOut4_47;
wire [7:0] nScanOut303;
wire [7:0] nOut4_48;
wire [7:0] nScanOut304;
wire [7:0] nOut4_49;
wire [7:0] nScanOut305;
wire [7:0] nOut4_50;
wire [7:0] nScanOut306;
wire [7:0] nOut4_51;
wire [7:0] nScanOut307;
wire [7:0] nOut4_52;
wire [7:0] nScanOut308;
wire [7:0] nOut4_53;
wire [7:0] nScanOut309;
wire [7:0] nOut4_54;
wire [7:0] nScanOut310;
wire [7:0] nOut4_55;
wire [7:0] nScanOut311;
wire [7:0] nOut4_56;
wire [7:0] nScanOut312;
wire [7:0] nOut4_57;
wire [7:0] nScanOut313;
wire [7:0] nOut4_58;
wire [7:0] nScanOut314;
wire [7:0] nOut4_59;
wire [7:0] nScanOut315;
wire [7:0] nOut4_60;
wire [7:0] nScanOut316;
wire [7:0] nOut4_61;
wire [7:0] nScanOut317;
wire [7:0] nOut4_62;
wire [7:0] nScanOut318;
wire [7:0] nOut4_63;
wire [7:0] nScanOut319;
wire [7:0] nOut5_0;
wire [7:0] nScanOut320;
wire [7:0] nOut5_1;
wire [7:0] nScanOut321;
wire [7:0] nOut5_2;
wire [7:0] nScanOut322;
wire [7:0] nOut5_3;
wire [7:0] nScanOut323;
wire [7:0] nOut5_4;
wire [7:0] nScanOut324;
wire [7:0] nOut5_5;
wire [7:0] nScanOut325;
wire [7:0] nOut5_6;
wire [7:0] nScanOut326;
wire [7:0] nOut5_7;
wire [7:0] nScanOut327;
wire [7:0] nOut5_8;
wire [7:0] nScanOut328;
wire [7:0] nOut5_9;
wire [7:0] nScanOut329;
wire [7:0] nOut5_10;
wire [7:0] nScanOut330;
wire [7:0] nOut5_11;
wire [7:0] nScanOut331;
wire [7:0] nOut5_12;
wire [7:0] nScanOut332;
wire [7:0] nOut5_13;
wire [7:0] nScanOut333;
wire [7:0] nOut5_14;
wire [7:0] nScanOut334;
wire [7:0] nOut5_15;
wire [7:0] nScanOut335;
wire [7:0] nOut5_16;
wire [7:0] nScanOut336;
wire [7:0] nOut5_17;
wire [7:0] nScanOut337;
wire [7:0] nOut5_18;
wire [7:0] nScanOut338;
wire [7:0] nOut5_19;
wire [7:0] nScanOut339;
wire [7:0] nOut5_20;
wire [7:0] nScanOut340;
wire [7:0] nOut5_21;
wire [7:0] nScanOut341;
wire [7:0] nOut5_22;
wire [7:0] nScanOut342;
wire [7:0] nOut5_23;
wire [7:0] nScanOut343;
wire [7:0] nOut5_24;
wire [7:0] nScanOut344;
wire [7:0] nOut5_25;
wire [7:0] nScanOut345;
wire [7:0] nOut5_26;
wire [7:0] nScanOut346;
wire [7:0] nOut5_27;
wire [7:0] nScanOut347;
wire [7:0] nOut5_28;
wire [7:0] nScanOut348;
wire [7:0] nOut5_29;
wire [7:0] nScanOut349;
wire [7:0] nOut5_30;
wire [7:0] nScanOut350;
wire [7:0] nOut5_31;
wire [7:0] nScanOut351;
wire [7:0] nOut5_32;
wire [7:0] nScanOut352;
wire [7:0] nOut5_33;
wire [7:0] nScanOut353;
wire [7:0] nOut5_34;
wire [7:0] nScanOut354;
wire [7:0] nOut5_35;
wire [7:0] nScanOut355;
wire [7:0] nOut5_36;
wire [7:0] nScanOut356;
wire [7:0] nOut5_37;
wire [7:0] nScanOut357;
wire [7:0] nOut5_38;
wire [7:0] nScanOut358;
wire [7:0] nOut5_39;
wire [7:0] nScanOut359;
wire [7:0] nOut5_40;
wire [7:0] nScanOut360;
wire [7:0] nOut5_41;
wire [7:0] nScanOut361;
wire [7:0] nOut5_42;
wire [7:0] nScanOut362;
wire [7:0] nOut5_43;
wire [7:0] nScanOut363;
wire [7:0] nOut5_44;
wire [7:0] nScanOut364;
wire [7:0] nOut5_45;
wire [7:0] nScanOut365;
wire [7:0] nOut5_46;
wire [7:0] nScanOut366;
wire [7:0] nOut5_47;
wire [7:0] nScanOut367;
wire [7:0] nOut5_48;
wire [7:0] nScanOut368;
wire [7:0] nOut5_49;
wire [7:0] nScanOut369;
wire [7:0] nOut5_50;
wire [7:0] nScanOut370;
wire [7:0] nOut5_51;
wire [7:0] nScanOut371;
wire [7:0] nOut5_52;
wire [7:0] nScanOut372;
wire [7:0] nOut5_53;
wire [7:0] nScanOut373;
wire [7:0] nOut5_54;
wire [7:0] nScanOut374;
wire [7:0] nOut5_55;
wire [7:0] nScanOut375;
wire [7:0] nOut5_56;
wire [7:0] nScanOut376;
wire [7:0] nOut5_57;
wire [7:0] nScanOut377;
wire [7:0] nOut5_58;
wire [7:0] nScanOut378;
wire [7:0] nOut5_59;
wire [7:0] nScanOut379;
wire [7:0] nOut5_60;
wire [7:0] nScanOut380;
wire [7:0] nOut5_61;
wire [7:0] nScanOut381;
wire [7:0] nOut5_62;
wire [7:0] nScanOut382;
wire [7:0] nOut5_63;
wire [7:0] nScanOut383;
wire [7:0] nOut6_0;
wire [7:0] nScanOut384;
wire [7:0] nOut6_1;
wire [7:0] nScanOut385;
wire [7:0] nOut6_2;
wire [7:0] nScanOut386;
wire [7:0] nOut6_3;
wire [7:0] nScanOut387;
wire [7:0] nOut6_4;
wire [7:0] nScanOut388;
wire [7:0] nOut6_5;
wire [7:0] nScanOut389;
wire [7:0] nOut6_6;
wire [7:0] nScanOut390;
wire [7:0] nOut6_7;
wire [7:0] nScanOut391;
wire [7:0] nOut6_8;
wire [7:0] nScanOut392;
wire [7:0] nOut6_9;
wire [7:0] nScanOut393;
wire [7:0] nOut6_10;
wire [7:0] nScanOut394;
wire [7:0] nOut6_11;
wire [7:0] nScanOut395;
wire [7:0] nOut6_12;
wire [7:0] nScanOut396;
wire [7:0] nOut6_13;
wire [7:0] nScanOut397;
wire [7:0] nOut6_14;
wire [7:0] nScanOut398;
wire [7:0] nOut6_15;
wire [7:0] nScanOut399;
wire [7:0] nOut6_16;
wire [7:0] nScanOut400;
wire [7:0] nOut6_17;
wire [7:0] nScanOut401;
wire [7:0] nOut6_18;
wire [7:0] nScanOut402;
wire [7:0] nOut6_19;
wire [7:0] nScanOut403;
wire [7:0] nOut6_20;
wire [7:0] nScanOut404;
wire [7:0] nOut6_21;
wire [7:0] nScanOut405;
wire [7:0] nOut6_22;
wire [7:0] nScanOut406;
wire [7:0] nOut6_23;
wire [7:0] nScanOut407;
wire [7:0] nOut6_24;
wire [7:0] nScanOut408;
wire [7:0] nOut6_25;
wire [7:0] nScanOut409;
wire [7:0] nOut6_26;
wire [7:0] nScanOut410;
wire [7:0] nOut6_27;
wire [7:0] nScanOut411;
wire [7:0] nOut6_28;
wire [7:0] nScanOut412;
wire [7:0] nOut6_29;
wire [7:0] nScanOut413;
wire [7:0] nOut6_30;
wire [7:0] nScanOut414;
wire [7:0] nOut6_31;
wire [7:0] nScanOut415;
wire [7:0] nOut6_32;
wire [7:0] nScanOut416;
wire [7:0] nOut6_33;
wire [7:0] nScanOut417;
wire [7:0] nOut6_34;
wire [7:0] nScanOut418;
wire [7:0] nOut6_35;
wire [7:0] nScanOut419;
wire [7:0] nOut6_36;
wire [7:0] nScanOut420;
wire [7:0] nOut6_37;
wire [7:0] nScanOut421;
wire [7:0] nOut6_38;
wire [7:0] nScanOut422;
wire [7:0] nOut6_39;
wire [7:0] nScanOut423;
wire [7:0] nOut6_40;
wire [7:0] nScanOut424;
wire [7:0] nOut6_41;
wire [7:0] nScanOut425;
wire [7:0] nOut6_42;
wire [7:0] nScanOut426;
wire [7:0] nOut6_43;
wire [7:0] nScanOut427;
wire [7:0] nOut6_44;
wire [7:0] nScanOut428;
wire [7:0] nOut6_45;
wire [7:0] nScanOut429;
wire [7:0] nOut6_46;
wire [7:0] nScanOut430;
wire [7:0] nOut6_47;
wire [7:0] nScanOut431;
wire [7:0] nOut6_48;
wire [7:0] nScanOut432;
wire [7:0] nOut6_49;
wire [7:0] nScanOut433;
wire [7:0] nOut6_50;
wire [7:0] nScanOut434;
wire [7:0] nOut6_51;
wire [7:0] nScanOut435;
wire [7:0] nOut6_52;
wire [7:0] nScanOut436;
wire [7:0] nOut6_53;
wire [7:0] nScanOut437;
wire [7:0] nOut6_54;
wire [7:0] nScanOut438;
wire [7:0] nOut6_55;
wire [7:0] nScanOut439;
wire [7:0] nOut6_56;
wire [7:0] nScanOut440;
wire [7:0] nOut6_57;
wire [7:0] nScanOut441;
wire [7:0] nOut6_58;
wire [7:0] nScanOut442;
wire [7:0] nOut6_59;
wire [7:0] nScanOut443;
wire [7:0] nOut6_60;
wire [7:0] nScanOut444;
wire [7:0] nOut6_61;
wire [7:0] nScanOut445;
wire [7:0] nOut6_62;
wire [7:0] nScanOut446;
wire [7:0] nOut6_63;
wire [7:0] nScanOut447;
wire [7:0] nOut7_0;
wire [7:0] nScanOut448;
wire [7:0] nOut7_1;
wire [7:0] nScanOut449;
wire [7:0] nOut7_2;
wire [7:0] nScanOut450;
wire [7:0] nOut7_3;
wire [7:0] nScanOut451;
wire [7:0] nOut7_4;
wire [7:0] nScanOut452;
wire [7:0] nOut7_5;
wire [7:0] nScanOut453;
wire [7:0] nOut7_6;
wire [7:0] nScanOut454;
wire [7:0] nOut7_7;
wire [7:0] nScanOut455;
wire [7:0] nOut7_8;
wire [7:0] nScanOut456;
wire [7:0] nOut7_9;
wire [7:0] nScanOut457;
wire [7:0] nOut7_10;
wire [7:0] nScanOut458;
wire [7:0] nOut7_11;
wire [7:0] nScanOut459;
wire [7:0] nOut7_12;
wire [7:0] nScanOut460;
wire [7:0] nOut7_13;
wire [7:0] nScanOut461;
wire [7:0] nOut7_14;
wire [7:0] nScanOut462;
wire [7:0] nOut7_15;
wire [7:0] nScanOut463;
wire [7:0] nOut7_16;
wire [7:0] nScanOut464;
wire [7:0] nOut7_17;
wire [7:0] nScanOut465;
wire [7:0] nOut7_18;
wire [7:0] nScanOut466;
wire [7:0] nOut7_19;
wire [7:0] nScanOut467;
wire [7:0] nOut7_20;
wire [7:0] nScanOut468;
wire [7:0] nOut7_21;
wire [7:0] nScanOut469;
wire [7:0] nOut7_22;
wire [7:0] nScanOut470;
wire [7:0] nOut7_23;
wire [7:0] nScanOut471;
wire [7:0] nOut7_24;
wire [7:0] nScanOut472;
wire [7:0] nOut7_25;
wire [7:0] nScanOut473;
wire [7:0] nOut7_26;
wire [7:0] nScanOut474;
wire [7:0] nOut7_27;
wire [7:0] nScanOut475;
wire [7:0] nOut7_28;
wire [7:0] nScanOut476;
wire [7:0] nOut7_29;
wire [7:0] nScanOut477;
wire [7:0] nOut7_30;
wire [7:0] nScanOut478;
wire [7:0] nOut7_31;
wire [7:0] nScanOut479;
wire [7:0] nOut7_32;
wire [7:0] nScanOut480;
wire [7:0] nOut7_33;
wire [7:0] nScanOut481;
wire [7:0] nOut7_34;
wire [7:0] nScanOut482;
wire [7:0] nOut7_35;
wire [7:0] nScanOut483;
wire [7:0] nOut7_36;
wire [7:0] nScanOut484;
wire [7:0] nOut7_37;
wire [7:0] nScanOut485;
wire [7:0] nOut7_38;
wire [7:0] nScanOut486;
wire [7:0] nOut7_39;
wire [7:0] nScanOut487;
wire [7:0] nOut7_40;
wire [7:0] nScanOut488;
wire [7:0] nOut7_41;
wire [7:0] nScanOut489;
wire [7:0] nOut7_42;
wire [7:0] nScanOut490;
wire [7:0] nOut7_43;
wire [7:0] nScanOut491;
wire [7:0] nOut7_44;
wire [7:0] nScanOut492;
wire [7:0] nOut7_45;
wire [7:0] nScanOut493;
wire [7:0] nOut7_46;
wire [7:0] nScanOut494;
wire [7:0] nOut7_47;
wire [7:0] nScanOut495;
wire [7:0] nOut7_48;
wire [7:0] nScanOut496;
wire [7:0] nOut7_49;
wire [7:0] nScanOut497;
wire [7:0] nOut7_50;
wire [7:0] nScanOut498;
wire [7:0] nOut7_51;
wire [7:0] nScanOut499;
wire [7:0] nOut7_52;
wire [7:0] nScanOut500;
wire [7:0] nOut7_53;
wire [7:0] nScanOut501;
wire [7:0] nOut7_54;
wire [7:0] nScanOut502;
wire [7:0] nOut7_55;
wire [7:0] nScanOut503;
wire [7:0] nOut7_56;
wire [7:0] nScanOut504;
wire [7:0] nOut7_57;
wire [7:0] nScanOut505;
wire [7:0] nOut7_58;
wire [7:0] nScanOut506;
wire [7:0] nOut7_59;
wire [7:0] nScanOut507;
wire [7:0] nOut7_60;
wire [7:0] nScanOut508;
wire [7:0] nOut7_61;
wire [7:0] nScanOut509;
wire [7:0] nOut7_62;
wire [7:0] nScanOut510;
wire [7:0] nOut7_63;
wire [7:0] nScanOut511;
wire [7:0] nOut8_0;
wire [7:0] nScanOut512;
wire [7:0] nOut8_1;
wire [7:0] nScanOut513;
wire [7:0] nOut8_2;
wire [7:0] nScanOut514;
wire [7:0] nOut8_3;
wire [7:0] nScanOut515;
wire [7:0] nOut8_4;
wire [7:0] nScanOut516;
wire [7:0] nOut8_5;
wire [7:0] nScanOut517;
wire [7:0] nOut8_6;
wire [7:0] nScanOut518;
wire [7:0] nOut8_7;
wire [7:0] nScanOut519;
wire [7:0] nOut8_8;
wire [7:0] nScanOut520;
wire [7:0] nOut8_9;
wire [7:0] nScanOut521;
wire [7:0] nOut8_10;
wire [7:0] nScanOut522;
wire [7:0] nOut8_11;
wire [7:0] nScanOut523;
wire [7:0] nOut8_12;
wire [7:0] nScanOut524;
wire [7:0] nOut8_13;
wire [7:0] nScanOut525;
wire [7:0] nOut8_14;
wire [7:0] nScanOut526;
wire [7:0] nOut8_15;
wire [7:0] nScanOut527;
wire [7:0] nOut8_16;
wire [7:0] nScanOut528;
wire [7:0] nOut8_17;
wire [7:0] nScanOut529;
wire [7:0] nOut8_18;
wire [7:0] nScanOut530;
wire [7:0] nOut8_19;
wire [7:0] nScanOut531;
wire [7:0] nOut8_20;
wire [7:0] nScanOut532;
wire [7:0] nOut8_21;
wire [7:0] nScanOut533;
wire [7:0] nOut8_22;
wire [7:0] nScanOut534;
wire [7:0] nOut8_23;
wire [7:0] nScanOut535;
wire [7:0] nOut8_24;
wire [7:0] nScanOut536;
wire [7:0] nOut8_25;
wire [7:0] nScanOut537;
wire [7:0] nOut8_26;
wire [7:0] nScanOut538;
wire [7:0] nOut8_27;
wire [7:0] nScanOut539;
wire [7:0] nOut8_28;
wire [7:0] nScanOut540;
wire [7:0] nOut8_29;
wire [7:0] nScanOut541;
wire [7:0] nOut8_30;
wire [7:0] nScanOut542;
wire [7:0] nOut8_31;
wire [7:0] nScanOut543;
wire [7:0] nOut8_32;
wire [7:0] nScanOut544;
wire [7:0] nOut8_33;
wire [7:0] nScanOut545;
wire [7:0] nOut8_34;
wire [7:0] nScanOut546;
wire [7:0] nOut8_35;
wire [7:0] nScanOut547;
wire [7:0] nOut8_36;
wire [7:0] nScanOut548;
wire [7:0] nOut8_37;
wire [7:0] nScanOut549;
wire [7:0] nOut8_38;
wire [7:0] nScanOut550;
wire [7:0] nOut8_39;
wire [7:0] nScanOut551;
wire [7:0] nOut8_40;
wire [7:0] nScanOut552;
wire [7:0] nOut8_41;
wire [7:0] nScanOut553;
wire [7:0] nOut8_42;
wire [7:0] nScanOut554;
wire [7:0] nOut8_43;
wire [7:0] nScanOut555;
wire [7:0] nOut8_44;
wire [7:0] nScanOut556;
wire [7:0] nOut8_45;
wire [7:0] nScanOut557;
wire [7:0] nOut8_46;
wire [7:0] nScanOut558;
wire [7:0] nOut8_47;
wire [7:0] nScanOut559;
wire [7:0] nOut8_48;
wire [7:0] nScanOut560;
wire [7:0] nOut8_49;
wire [7:0] nScanOut561;
wire [7:0] nOut8_50;
wire [7:0] nScanOut562;
wire [7:0] nOut8_51;
wire [7:0] nScanOut563;
wire [7:0] nOut8_52;
wire [7:0] nScanOut564;
wire [7:0] nOut8_53;
wire [7:0] nScanOut565;
wire [7:0] nOut8_54;
wire [7:0] nScanOut566;
wire [7:0] nOut8_55;
wire [7:0] nScanOut567;
wire [7:0] nOut8_56;
wire [7:0] nScanOut568;
wire [7:0] nOut8_57;
wire [7:0] nScanOut569;
wire [7:0] nOut8_58;
wire [7:0] nScanOut570;
wire [7:0] nOut8_59;
wire [7:0] nScanOut571;
wire [7:0] nOut8_60;
wire [7:0] nScanOut572;
wire [7:0] nOut8_61;
wire [7:0] nScanOut573;
wire [7:0] nOut8_62;
wire [7:0] nScanOut574;
wire [7:0] nOut8_63;
wire [7:0] nScanOut575;
wire [7:0] nOut9_0;
wire [7:0] nScanOut576;
wire [7:0] nOut9_1;
wire [7:0] nScanOut577;
wire [7:0] nOut9_2;
wire [7:0] nScanOut578;
wire [7:0] nOut9_3;
wire [7:0] nScanOut579;
wire [7:0] nOut9_4;
wire [7:0] nScanOut580;
wire [7:0] nOut9_5;
wire [7:0] nScanOut581;
wire [7:0] nOut9_6;
wire [7:0] nScanOut582;
wire [7:0] nOut9_7;
wire [7:0] nScanOut583;
wire [7:0] nOut9_8;
wire [7:0] nScanOut584;
wire [7:0] nOut9_9;
wire [7:0] nScanOut585;
wire [7:0] nOut9_10;
wire [7:0] nScanOut586;
wire [7:0] nOut9_11;
wire [7:0] nScanOut587;
wire [7:0] nOut9_12;
wire [7:0] nScanOut588;
wire [7:0] nOut9_13;
wire [7:0] nScanOut589;
wire [7:0] nOut9_14;
wire [7:0] nScanOut590;
wire [7:0] nOut9_15;
wire [7:0] nScanOut591;
wire [7:0] nOut9_16;
wire [7:0] nScanOut592;
wire [7:0] nOut9_17;
wire [7:0] nScanOut593;
wire [7:0] nOut9_18;
wire [7:0] nScanOut594;
wire [7:0] nOut9_19;
wire [7:0] nScanOut595;
wire [7:0] nOut9_20;
wire [7:0] nScanOut596;
wire [7:0] nOut9_21;
wire [7:0] nScanOut597;
wire [7:0] nOut9_22;
wire [7:0] nScanOut598;
wire [7:0] nOut9_23;
wire [7:0] nScanOut599;
wire [7:0] nOut9_24;
wire [7:0] nScanOut600;
wire [7:0] nOut9_25;
wire [7:0] nScanOut601;
wire [7:0] nOut9_26;
wire [7:0] nScanOut602;
wire [7:0] nOut9_27;
wire [7:0] nScanOut603;
wire [7:0] nOut9_28;
wire [7:0] nScanOut604;
wire [7:0] nOut9_29;
wire [7:0] nScanOut605;
wire [7:0] nOut9_30;
wire [7:0] nScanOut606;
wire [7:0] nOut9_31;
wire [7:0] nScanOut607;
wire [7:0] nOut9_32;
wire [7:0] nScanOut608;
wire [7:0] nOut9_33;
wire [7:0] nScanOut609;
wire [7:0] nOut9_34;
wire [7:0] nScanOut610;
wire [7:0] nOut9_35;
wire [7:0] nScanOut611;
wire [7:0] nOut9_36;
wire [7:0] nScanOut612;
wire [7:0] nOut9_37;
wire [7:0] nScanOut613;
wire [7:0] nOut9_38;
wire [7:0] nScanOut614;
wire [7:0] nOut9_39;
wire [7:0] nScanOut615;
wire [7:0] nOut9_40;
wire [7:0] nScanOut616;
wire [7:0] nOut9_41;
wire [7:0] nScanOut617;
wire [7:0] nOut9_42;
wire [7:0] nScanOut618;
wire [7:0] nOut9_43;
wire [7:0] nScanOut619;
wire [7:0] nOut9_44;
wire [7:0] nScanOut620;
wire [7:0] nOut9_45;
wire [7:0] nScanOut621;
wire [7:0] nOut9_46;
wire [7:0] nScanOut622;
wire [7:0] nOut9_47;
wire [7:0] nScanOut623;
wire [7:0] nOut9_48;
wire [7:0] nScanOut624;
wire [7:0] nOut9_49;
wire [7:0] nScanOut625;
wire [7:0] nOut9_50;
wire [7:0] nScanOut626;
wire [7:0] nOut9_51;
wire [7:0] nScanOut627;
wire [7:0] nOut9_52;
wire [7:0] nScanOut628;
wire [7:0] nOut9_53;
wire [7:0] nScanOut629;
wire [7:0] nOut9_54;
wire [7:0] nScanOut630;
wire [7:0] nOut9_55;
wire [7:0] nScanOut631;
wire [7:0] nOut9_56;
wire [7:0] nScanOut632;
wire [7:0] nOut9_57;
wire [7:0] nScanOut633;
wire [7:0] nOut9_58;
wire [7:0] nScanOut634;
wire [7:0] nOut9_59;
wire [7:0] nScanOut635;
wire [7:0] nOut9_60;
wire [7:0] nScanOut636;
wire [7:0] nOut9_61;
wire [7:0] nScanOut637;
wire [7:0] nOut9_62;
wire [7:0] nScanOut638;
wire [7:0] nOut9_63;
wire [7:0] nScanOut639;
wire [7:0] nOut10_0;
wire [7:0] nScanOut640;
wire [7:0] nOut10_1;
wire [7:0] nScanOut641;
wire [7:0] nOut10_2;
wire [7:0] nScanOut642;
wire [7:0] nOut10_3;
wire [7:0] nScanOut643;
wire [7:0] nOut10_4;
wire [7:0] nScanOut644;
wire [7:0] nOut10_5;
wire [7:0] nScanOut645;
wire [7:0] nOut10_6;
wire [7:0] nScanOut646;
wire [7:0] nOut10_7;
wire [7:0] nScanOut647;
wire [7:0] nOut10_8;
wire [7:0] nScanOut648;
wire [7:0] nOut10_9;
wire [7:0] nScanOut649;
wire [7:0] nOut10_10;
wire [7:0] nScanOut650;
wire [7:0] nOut10_11;
wire [7:0] nScanOut651;
wire [7:0] nOut10_12;
wire [7:0] nScanOut652;
wire [7:0] nOut10_13;
wire [7:0] nScanOut653;
wire [7:0] nOut10_14;
wire [7:0] nScanOut654;
wire [7:0] nOut10_15;
wire [7:0] nScanOut655;
wire [7:0] nOut10_16;
wire [7:0] nScanOut656;
wire [7:0] nOut10_17;
wire [7:0] nScanOut657;
wire [7:0] nOut10_18;
wire [7:0] nScanOut658;
wire [7:0] nOut10_19;
wire [7:0] nScanOut659;
wire [7:0] nOut10_20;
wire [7:0] nScanOut660;
wire [7:0] nOut10_21;
wire [7:0] nScanOut661;
wire [7:0] nOut10_22;
wire [7:0] nScanOut662;
wire [7:0] nOut10_23;
wire [7:0] nScanOut663;
wire [7:0] nOut10_24;
wire [7:0] nScanOut664;
wire [7:0] nOut10_25;
wire [7:0] nScanOut665;
wire [7:0] nOut10_26;
wire [7:0] nScanOut666;
wire [7:0] nOut10_27;
wire [7:0] nScanOut667;
wire [7:0] nOut10_28;
wire [7:0] nScanOut668;
wire [7:0] nOut10_29;
wire [7:0] nScanOut669;
wire [7:0] nOut10_30;
wire [7:0] nScanOut670;
wire [7:0] nOut10_31;
wire [7:0] nScanOut671;
wire [7:0] nOut10_32;
wire [7:0] nScanOut672;
wire [7:0] nOut10_33;
wire [7:0] nScanOut673;
wire [7:0] nOut10_34;
wire [7:0] nScanOut674;
wire [7:0] nOut10_35;
wire [7:0] nScanOut675;
wire [7:0] nOut10_36;
wire [7:0] nScanOut676;
wire [7:0] nOut10_37;
wire [7:0] nScanOut677;
wire [7:0] nOut10_38;
wire [7:0] nScanOut678;
wire [7:0] nOut10_39;
wire [7:0] nScanOut679;
wire [7:0] nOut10_40;
wire [7:0] nScanOut680;
wire [7:0] nOut10_41;
wire [7:0] nScanOut681;
wire [7:0] nOut10_42;
wire [7:0] nScanOut682;
wire [7:0] nOut10_43;
wire [7:0] nScanOut683;
wire [7:0] nOut10_44;
wire [7:0] nScanOut684;
wire [7:0] nOut10_45;
wire [7:0] nScanOut685;
wire [7:0] nOut10_46;
wire [7:0] nScanOut686;
wire [7:0] nOut10_47;
wire [7:0] nScanOut687;
wire [7:0] nOut10_48;
wire [7:0] nScanOut688;
wire [7:0] nOut10_49;
wire [7:0] nScanOut689;
wire [7:0] nOut10_50;
wire [7:0] nScanOut690;
wire [7:0] nOut10_51;
wire [7:0] nScanOut691;
wire [7:0] nOut10_52;
wire [7:0] nScanOut692;
wire [7:0] nOut10_53;
wire [7:0] nScanOut693;
wire [7:0] nOut10_54;
wire [7:0] nScanOut694;
wire [7:0] nOut10_55;
wire [7:0] nScanOut695;
wire [7:0] nOut10_56;
wire [7:0] nScanOut696;
wire [7:0] nOut10_57;
wire [7:0] nScanOut697;
wire [7:0] nOut10_58;
wire [7:0] nScanOut698;
wire [7:0] nOut10_59;
wire [7:0] nScanOut699;
wire [7:0] nOut10_60;
wire [7:0] nScanOut700;
wire [7:0] nOut10_61;
wire [7:0] nScanOut701;
wire [7:0] nOut10_62;
wire [7:0] nScanOut702;
wire [7:0] nOut10_63;
wire [7:0] nScanOut703;
wire [7:0] nOut11_0;
wire [7:0] nScanOut704;
wire [7:0] nOut11_1;
wire [7:0] nScanOut705;
wire [7:0] nOut11_2;
wire [7:0] nScanOut706;
wire [7:0] nOut11_3;
wire [7:0] nScanOut707;
wire [7:0] nOut11_4;
wire [7:0] nScanOut708;
wire [7:0] nOut11_5;
wire [7:0] nScanOut709;
wire [7:0] nOut11_6;
wire [7:0] nScanOut710;
wire [7:0] nOut11_7;
wire [7:0] nScanOut711;
wire [7:0] nOut11_8;
wire [7:0] nScanOut712;
wire [7:0] nOut11_9;
wire [7:0] nScanOut713;
wire [7:0] nOut11_10;
wire [7:0] nScanOut714;
wire [7:0] nOut11_11;
wire [7:0] nScanOut715;
wire [7:0] nOut11_12;
wire [7:0] nScanOut716;
wire [7:0] nOut11_13;
wire [7:0] nScanOut717;
wire [7:0] nOut11_14;
wire [7:0] nScanOut718;
wire [7:0] nOut11_15;
wire [7:0] nScanOut719;
wire [7:0] nOut11_16;
wire [7:0] nScanOut720;
wire [7:0] nOut11_17;
wire [7:0] nScanOut721;
wire [7:0] nOut11_18;
wire [7:0] nScanOut722;
wire [7:0] nOut11_19;
wire [7:0] nScanOut723;
wire [7:0] nOut11_20;
wire [7:0] nScanOut724;
wire [7:0] nOut11_21;
wire [7:0] nScanOut725;
wire [7:0] nOut11_22;
wire [7:0] nScanOut726;
wire [7:0] nOut11_23;
wire [7:0] nScanOut727;
wire [7:0] nOut11_24;
wire [7:0] nScanOut728;
wire [7:0] nOut11_25;
wire [7:0] nScanOut729;
wire [7:0] nOut11_26;
wire [7:0] nScanOut730;
wire [7:0] nOut11_27;
wire [7:0] nScanOut731;
wire [7:0] nOut11_28;
wire [7:0] nScanOut732;
wire [7:0] nOut11_29;
wire [7:0] nScanOut733;
wire [7:0] nOut11_30;
wire [7:0] nScanOut734;
wire [7:0] nOut11_31;
wire [7:0] nScanOut735;
wire [7:0] nOut11_32;
wire [7:0] nScanOut736;
wire [7:0] nOut11_33;
wire [7:0] nScanOut737;
wire [7:0] nOut11_34;
wire [7:0] nScanOut738;
wire [7:0] nOut11_35;
wire [7:0] nScanOut739;
wire [7:0] nOut11_36;
wire [7:0] nScanOut740;
wire [7:0] nOut11_37;
wire [7:0] nScanOut741;
wire [7:0] nOut11_38;
wire [7:0] nScanOut742;
wire [7:0] nOut11_39;
wire [7:0] nScanOut743;
wire [7:0] nOut11_40;
wire [7:0] nScanOut744;
wire [7:0] nOut11_41;
wire [7:0] nScanOut745;
wire [7:0] nOut11_42;
wire [7:0] nScanOut746;
wire [7:0] nOut11_43;
wire [7:0] nScanOut747;
wire [7:0] nOut11_44;
wire [7:0] nScanOut748;
wire [7:0] nOut11_45;
wire [7:0] nScanOut749;
wire [7:0] nOut11_46;
wire [7:0] nScanOut750;
wire [7:0] nOut11_47;
wire [7:0] nScanOut751;
wire [7:0] nOut11_48;
wire [7:0] nScanOut752;
wire [7:0] nOut11_49;
wire [7:0] nScanOut753;
wire [7:0] nOut11_50;
wire [7:0] nScanOut754;
wire [7:0] nOut11_51;
wire [7:0] nScanOut755;
wire [7:0] nOut11_52;
wire [7:0] nScanOut756;
wire [7:0] nOut11_53;
wire [7:0] nScanOut757;
wire [7:0] nOut11_54;
wire [7:0] nScanOut758;
wire [7:0] nOut11_55;
wire [7:0] nScanOut759;
wire [7:0] nOut11_56;
wire [7:0] nScanOut760;
wire [7:0] nOut11_57;
wire [7:0] nScanOut761;
wire [7:0] nOut11_58;
wire [7:0] nScanOut762;
wire [7:0] nOut11_59;
wire [7:0] nScanOut763;
wire [7:0] nOut11_60;
wire [7:0] nScanOut764;
wire [7:0] nOut11_61;
wire [7:0] nScanOut765;
wire [7:0] nOut11_62;
wire [7:0] nScanOut766;
wire [7:0] nOut11_63;
wire [7:0] nScanOut767;
wire [7:0] nOut12_0;
wire [7:0] nScanOut768;
wire [7:0] nOut12_1;
wire [7:0] nScanOut769;
wire [7:0] nOut12_2;
wire [7:0] nScanOut770;
wire [7:0] nOut12_3;
wire [7:0] nScanOut771;
wire [7:0] nOut12_4;
wire [7:0] nScanOut772;
wire [7:0] nOut12_5;
wire [7:0] nScanOut773;
wire [7:0] nOut12_6;
wire [7:0] nScanOut774;
wire [7:0] nOut12_7;
wire [7:0] nScanOut775;
wire [7:0] nOut12_8;
wire [7:0] nScanOut776;
wire [7:0] nOut12_9;
wire [7:0] nScanOut777;
wire [7:0] nOut12_10;
wire [7:0] nScanOut778;
wire [7:0] nOut12_11;
wire [7:0] nScanOut779;
wire [7:0] nOut12_12;
wire [7:0] nScanOut780;
wire [7:0] nOut12_13;
wire [7:0] nScanOut781;
wire [7:0] nOut12_14;
wire [7:0] nScanOut782;
wire [7:0] nOut12_15;
wire [7:0] nScanOut783;
wire [7:0] nOut12_16;
wire [7:0] nScanOut784;
wire [7:0] nOut12_17;
wire [7:0] nScanOut785;
wire [7:0] nOut12_18;
wire [7:0] nScanOut786;
wire [7:0] nOut12_19;
wire [7:0] nScanOut787;
wire [7:0] nOut12_20;
wire [7:0] nScanOut788;
wire [7:0] nOut12_21;
wire [7:0] nScanOut789;
wire [7:0] nOut12_22;
wire [7:0] nScanOut790;
wire [7:0] nOut12_23;
wire [7:0] nScanOut791;
wire [7:0] nOut12_24;
wire [7:0] nScanOut792;
wire [7:0] nOut12_25;
wire [7:0] nScanOut793;
wire [7:0] nOut12_26;
wire [7:0] nScanOut794;
wire [7:0] nOut12_27;
wire [7:0] nScanOut795;
wire [7:0] nOut12_28;
wire [7:0] nScanOut796;
wire [7:0] nOut12_29;
wire [7:0] nScanOut797;
wire [7:0] nOut12_30;
wire [7:0] nScanOut798;
wire [7:0] nOut12_31;
wire [7:0] nScanOut799;
wire [7:0] nOut12_32;
wire [7:0] nScanOut800;
wire [7:0] nOut12_33;
wire [7:0] nScanOut801;
wire [7:0] nOut12_34;
wire [7:0] nScanOut802;
wire [7:0] nOut12_35;
wire [7:0] nScanOut803;
wire [7:0] nOut12_36;
wire [7:0] nScanOut804;
wire [7:0] nOut12_37;
wire [7:0] nScanOut805;
wire [7:0] nOut12_38;
wire [7:0] nScanOut806;
wire [7:0] nOut12_39;
wire [7:0] nScanOut807;
wire [7:0] nOut12_40;
wire [7:0] nScanOut808;
wire [7:0] nOut12_41;
wire [7:0] nScanOut809;
wire [7:0] nOut12_42;
wire [7:0] nScanOut810;
wire [7:0] nOut12_43;
wire [7:0] nScanOut811;
wire [7:0] nOut12_44;
wire [7:0] nScanOut812;
wire [7:0] nOut12_45;
wire [7:0] nScanOut813;
wire [7:0] nOut12_46;
wire [7:0] nScanOut814;
wire [7:0] nOut12_47;
wire [7:0] nScanOut815;
wire [7:0] nOut12_48;
wire [7:0] nScanOut816;
wire [7:0] nOut12_49;
wire [7:0] nScanOut817;
wire [7:0] nOut12_50;
wire [7:0] nScanOut818;
wire [7:0] nOut12_51;
wire [7:0] nScanOut819;
wire [7:0] nOut12_52;
wire [7:0] nScanOut820;
wire [7:0] nOut12_53;
wire [7:0] nScanOut821;
wire [7:0] nOut12_54;
wire [7:0] nScanOut822;
wire [7:0] nOut12_55;
wire [7:0] nScanOut823;
wire [7:0] nOut12_56;
wire [7:0] nScanOut824;
wire [7:0] nOut12_57;
wire [7:0] nScanOut825;
wire [7:0] nOut12_58;
wire [7:0] nScanOut826;
wire [7:0] nOut12_59;
wire [7:0] nScanOut827;
wire [7:0] nOut12_60;
wire [7:0] nScanOut828;
wire [7:0] nOut12_61;
wire [7:0] nScanOut829;
wire [7:0] nOut12_62;
wire [7:0] nScanOut830;
wire [7:0] nOut12_63;
wire [7:0] nScanOut831;
wire [7:0] nOut13_0;
wire [7:0] nScanOut832;
wire [7:0] nOut13_1;
wire [7:0] nScanOut833;
wire [7:0] nOut13_2;
wire [7:0] nScanOut834;
wire [7:0] nOut13_3;
wire [7:0] nScanOut835;
wire [7:0] nOut13_4;
wire [7:0] nScanOut836;
wire [7:0] nOut13_5;
wire [7:0] nScanOut837;
wire [7:0] nOut13_6;
wire [7:0] nScanOut838;
wire [7:0] nOut13_7;
wire [7:0] nScanOut839;
wire [7:0] nOut13_8;
wire [7:0] nScanOut840;
wire [7:0] nOut13_9;
wire [7:0] nScanOut841;
wire [7:0] nOut13_10;
wire [7:0] nScanOut842;
wire [7:0] nOut13_11;
wire [7:0] nScanOut843;
wire [7:0] nOut13_12;
wire [7:0] nScanOut844;
wire [7:0] nOut13_13;
wire [7:0] nScanOut845;
wire [7:0] nOut13_14;
wire [7:0] nScanOut846;
wire [7:0] nOut13_15;
wire [7:0] nScanOut847;
wire [7:0] nOut13_16;
wire [7:0] nScanOut848;
wire [7:0] nOut13_17;
wire [7:0] nScanOut849;
wire [7:0] nOut13_18;
wire [7:0] nScanOut850;
wire [7:0] nOut13_19;
wire [7:0] nScanOut851;
wire [7:0] nOut13_20;
wire [7:0] nScanOut852;
wire [7:0] nOut13_21;
wire [7:0] nScanOut853;
wire [7:0] nOut13_22;
wire [7:0] nScanOut854;
wire [7:0] nOut13_23;
wire [7:0] nScanOut855;
wire [7:0] nOut13_24;
wire [7:0] nScanOut856;
wire [7:0] nOut13_25;
wire [7:0] nScanOut857;
wire [7:0] nOut13_26;
wire [7:0] nScanOut858;
wire [7:0] nOut13_27;
wire [7:0] nScanOut859;
wire [7:0] nOut13_28;
wire [7:0] nScanOut860;
wire [7:0] nOut13_29;
wire [7:0] nScanOut861;
wire [7:0] nOut13_30;
wire [7:0] nScanOut862;
wire [7:0] nOut13_31;
wire [7:0] nScanOut863;
wire [7:0] nOut13_32;
wire [7:0] nScanOut864;
wire [7:0] nOut13_33;
wire [7:0] nScanOut865;
wire [7:0] nOut13_34;
wire [7:0] nScanOut866;
wire [7:0] nOut13_35;
wire [7:0] nScanOut867;
wire [7:0] nOut13_36;
wire [7:0] nScanOut868;
wire [7:0] nOut13_37;
wire [7:0] nScanOut869;
wire [7:0] nOut13_38;
wire [7:0] nScanOut870;
wire [7:0] nOut13_39;
wire [7:0] nScanOut871;
wire [7:0] nOut13_40;
wire [7:0] nScanOut872;
wire [7:0] nOut13_41;
wire [7:0] nScanOut873;
wire [7:0] nOut13_42;
wire [7:0] nScanOut874;
wire [7:0] nOut13_43;
wire [7:0] nScanOut875;
wire [7:0] nOut13_44;
wire [7:0] nScanOut876;
wire [7:0] nOut13_45;
wire [7:0] nScanOut877;
wire [7:0] nOut13_46;
wire [7:0] nScanOut878;
wire [7:0] nOut13_47;
wire [7:0] nScanOut879;
wire [7:0] nOut13_48;
wire [7:0] nScanOut880;
wire [7:0] nOut13_49;
wire [7:0] nScanOut881;
wire [7:0] nOut13_50;
wire [7:0] nScanOut882;
wire [7:0] nOut13_51;
wire [7:0] nScanOut883;
wire [7:0] nOut13_52;
wire [7:0] nScanOut884;
wire [7:0] nOut13_53;
wire [7:0] nScanOut885;
wire [7:0] nOut13_54;
wire [7:0] nScanOut886;
wire [7:0] nOut13_55;
wire [7:0] nScanOut887;
wire [7:0] nOut13_56;
wire [7:0] nScanOut888;
wire [7:0] nOut13_57;
wire [7:0] nScanOut889;
wire [7:0] nOut13_58;
wire [7:0] nScanOut890;
wire [7:0] nOut13_59;
wire [7:0] nScanOut891;
wire [7:0] nOut13_60;
wire [7:0] nScanOut892;
wire [7:0] nOut13_61;
wire [7:0] nScanOut893;
wire [7:0] nOut13_62;
wire [7:0] nScanOut894;
wire [7:0] nOut13_63;
wire [7:0] nScanOut895;
wire [7:0] nOut14_0;
wire [7:0] nScanOut896;
wire [7:0] nOut14_1;
wire [7:0] nScanOut897;
wire [7:0] nOut14_2;
wire [7:0] nScanOut898;
wire [7:0] nOut14_3;
wire [7:0] nScanOut899;
wire [7:0] nOut14_4;
wire [7:0] nScanOut900;
wire [7:0] nOut14_5;
wire [7:0] nScanOut901;
wire [7:0] nOut14_6;
wire [7:0] nScanOut902;
wire [7:0] nOut14_7;
wire [7:0] nScanOut903;
wire [7:0] nOut14_8;
wire [7:0] nScanOut904;
wire [7:0] nOut14_9;
wire [7:0] nScanOut905;
wire [7:0] nOut14_10;
wire [7:0] nScanOut906;
wire [7:0] nOut14_11;
wire [7:0] nScanOut907;
wire [7:0] nOut14_12;
wire [7:0] nScanOut908;
wire [7:0] nOut14_13;
wire [7:0] nScanOut909;
wire [7:0] nOut14_14;
wire [7:0] nScanOut910;
wire [7:0] nOut14_15;
wire [7:0] nScanOut911;
wire [7:0] nOut14_16;
wire [7:0] nScanOut912;
wire [7:0] nOut14_17;
wire [7:0] nScanOut913;
wire [7:0] nOut14_18;
wire [7:0] nScanOut914;
wire [7:0] nOut14_19;
wire [7:0] nScanOut915;
wire [7:0] nOut14_20;
wire [7:0] nScanOut916;
wire [7:0] nOut14_21;
wire [7:0] nScanOut917;
wire [7:0] nOut14_22;
wire [7:0] nScanOut918;
wire [7:0] nOut14_23;
wire [7:0] nScanOut919;
wire [7:0] nOut14_24;
wire [7:0] nScanOut920;
wire [7:0] nOut14_25;
wire [7:0] nScanOut921;
wire [7:0] nOut14_26;
wire [7:0] nScanOut922;
wire [7:0] nOut14_27;
wire [7:0] nScanOut923;
wire [7:0] nOut14_28;
wire [7:0] nScanOut924;
wire [7:0] nOut14_29;
wire [7:0] nScanOut925;
wire [7:0] nOut14_30;
wire [7:0] nScanOut926;
wire [7:0] nOut14_31;
wire [7:0] nScanOut927;
wire [7:0] nOut14_32;
wire [7:0] nScanOut928;
wire [7:0] nOut14_33;
wire [7:0] nScanOut929;
wire [7:0] nOut14_34;
wire [7:0] nScanOut930;
wire [7:0] nOut14_35;
wire [7:0] nScanOut931;
wire [7:0] nOut14_36;
wire [7:0] nScanOut932;
wire [7:0] nOut14_37;
wire [7:0] nScanOut933;
wire [7:0] nOut14_38;
wire [7:0] nScanOut934;
wire [7:0] nOut14_39;
wire [7:0] nScanOut935;
wire [7:0] nOut14_40;
wire [7:0] nScanOut936;
wire [7:0] nOut14_41;
wire [7:0] nScanOut937;
wire [7:0] nOut14_42;
wire [7:0] nScanOut938;
wire [7:0] nOut14_43;
wire [7:0] nScanOut939;
wire [7:0] nOut14_44;
wire [7:0] nScanOut940;
wire [7:0] nOut14_45;
wire [7:0] nScanOut941;
wire [7:0] nOut14_46;
wire [7:0] nScanOut942;
wire [7:0] nOut14_47;
wire [7:0] nScanOut943;
wire [7:0] nOut14_48;
wire [7:0] nScanOut944;
wire [7:0] nOut14_49;
wire [7:0] nScanOut945;
wire [7:0] nOut14_50;
wire [7:0] nScanOut946;
wire [7:0] nOut14_51;
wire [7:0] nScanOut947;
wire [7:0] nOut14_52;
wire [7:0] nScanOut948;
wire [7:0] nOut14_53;
wire [7:0] nScanOut949;
wire [7:0] nOut14_54;
wire [7:0] nScanOut950;
wire [7:0] nOut14_55;
wire [7:0] nScanOut951;
wire [7:0] nOut14_56;
wire [7:0] nScanOut952;
wire [7:0] nOut14_57;
wire [7:0] nScanOut953;
wire [7:0] nOut14_58;
wire [7:0] nScanOut954;
wire [7:0] nOut14_59;
wire [7:0] nScanOut955;
wire [7:0] nOut14_60;
wire [7:0] nScanOut956;
wire [7:0] nOut14_61;
wire [7:0] nScanOut957;
wire [7:0] nOut14_62;
wire [7:0] nScanOut958;
wire [7:0] nOut14_63;
wire [7:0] nScanOut959;
wire [7:0] nOut15_0;
wire [7:0] nScanOut960;
wire [7:0] nOut15_1;
wire [7:0] nScanOut961;
wire [7:0] nOut15_2;
wire [7:0] nScanOut962;
wire [7:0] nOut15_3;
wire [7:0] nScanOut963;
wire [7:0] nOut15_4;
wire [7:0] nScanOut964;
wire [7:0] nOut15_5;
wire [7:0] nScanOut965;
wire [7:0] nOut15_6;
wire [7:0] nScanOut966;
wire [7:0] nOut15_7;
wire [7:0] nScanOut967;
wire [7:0] nOut15_8;
wire [7:0] nScanOut968;
wire [7:0] nOut15_9;
wire [7:0] nScanOut969;
wire [7:0] nOut15_10;
wire [7:0] nScanOut970;
wire [7:0] nOut15_11;
wire [7:0] nScanOut971;
wire [7:0] nOut15_12;
wire [7:0] nScanOut972;
wire [7:0] nOut15_13;
wire [7:0] nScanOut973;
wire [7:0] nOut15_14;
wire [7:0] nScanOut974;
wire [7:0] nOut15_15;
wire [7:0] nScanOut975;
wire [7:0] nOut15_16;
wire [7:0] nScanOut976;
wire [7:0] nOut15_17;
wire [7:0] nScanOut977;
wire [7:0] nOut15_18;
wire [7:0] nScanOut978;
wire [7:0] nOut15_19;
wire [7:0] nScanOut979;
wire [7:0] nOut15_20;
wire [7:0] nScanOut980;
wire [7:0] nOut15_21;
wire [7:0] nScanOut981;
wire [7:0] nOut15_22;
wire [7:0] nScanOut982;
wire [7:0] nOut15_23;
wire [7:0] nScanOut983;
wire [7:0] nOut15_24;
wire [7:0] nScanOut984;
wire [7:0] nOut15_25;
wire [7:0] nScanOut985;
wire [7:0] nOut15_26;
wire [7:0] nScanOut986;
wire [7:0] nOut15_27;
wire [7:0] nScanOut987;
wire [7:0] nOut15_28;
wire [7:0] nScanOut988;
wire [7:0] nOut15_29;
wire [7:0] nScanOut989;
wire [7:0] nOut15_30;
wire [7:0] nScanOut990;
wire [7:0] nOut15_31;
wire [7:0] nScanOut991;
wire [7:0] nOut15_32;
wire [7:0] nScanOut992;
wire [7:0] nOut15_33;
wire [7:0] nScanOut993;
wire [7:0] nOut15_34;
wire [7:0] nScanOut994;
wire [7:0] nOut15_35;
wire [7:0] nScanOut995;
wire [7:0] nOut15_36;
wire [7:0] nScanOut996;
wire [7:0] nOut15_37;
wire [7:0] nScanOut997;
wire [7:0] nOut15_38;
wire [7:0] nScanOut998;
wire [7:0] nOut15_39;
wire [7:0] nScanOut999;
wire [7:0] nOut15_40;
wire [7:0] nScanOut1000;
wire [7:0] nOut15_41;
wire [7:0] nScanOut1001;
wire [7:0] nOut15_42;
wire [7:0] nScanOut1002;
wire [7:0] nOut15_43;
wire [7:0] nScanOut1003;
wire [7:0] nOut15_44;
wire [7:0] nScanOut1004;
wire [7:0] nOut15_45;
wire [7:0] nScanOut1005;
wire [7:0] nOut15_46;
wire [7:0] nScanOut1006;
wire [7:0] nOut15_47;
wire [7:0] nScanOut1007;
wire [7:0] nOut15_48;
wire [7:0] nScanOut1008;
wire [7:0] nOut15_49;
wire [7:0] nScanOut1009;
wire [7:0] nOut15_50;
wire [7:0] nScanOut1010;
wire [7:0] nOut15_51;
wire [7:0] nScanOut1011;
wire [7:0] nOut15_52;
wire [7:0] nScanOut1012;
wire [7:0] nOut15_53;
wire [7:0] nScanOut1013;
wire [7:0] nOut15_54;
wire [7:0] nScanOut1014;
wire [7:0] nOut15_55;
wire [7:0] nScanOut1015;
wire [7:0] nOut15_56;
wire [7:0] nScanOut1016;
wire [7:0] nOut15_57;
wire [7:0] nScanOut1017;
wire [7:0] nOut15_58;
wire [7:0] nScanOut1018;
wire [7:0] nOut15_59;
wire [7:0] nScanOut1019;
wire [7:0] nOut15_60;
wire [7:0] nScanOut1020;
wire [7:0] nOut15_61;
wire [7:0] nScanOut1021;
wire [7:0] nOut15_62;
wire [7:0] nScanOut1022;
wire [7:0] nOut15_63;
wire [7:0] nScanOut1023;
wire [7:0] nOut16_0;
wire [7:0] nScanOut1024;
wire [7:0] nOut16_1;
wire [7:0] nScanOut1025;
wire [7:0] nOut16_2;
wire [7:0] nScanOut1026;
wire [7:0] nOut16_3;
wire [7:0] nScanOut1027;
wire [7:0] nOut16_4;
wire [7:0] nScanOut1028;
wire [7:0] nOut16_5;
wire [7:0] nScanOut1029;
wire [7:0] nOut16_6;
wire [7:0] nScanOut1030;
wire [7:0] nOut16_7;
wire [7:0] nScanOut1031;
wire [7:0] nOut16_8;
wire [7:0] nScanOut1032;
wire [7:0] nOut16_9;
wire [7:0] nScanOut1033;
wire [7:0] nOut16_10;
wire [7:0] nScanOut1034;
wire [7:0] nOut16_11;
wire [7:0] nScanOut1035;
wire [7:0] nOut16_12;
wire [7:0] nScanOut1036;
wire [7:0] nOut16_13;
wire [7:0] nScanOut1037;
wire [7:0] nOut16_14;
wire [7:0] nScanOut1038;
wire [7:0] nOut16_15;
wire [7:0] nScanOut1039;
wire [7:0] nOut16_16;
wire [7:0] nScanOut1040;
wire [7:0] nOut16_17;
wire [7:0] nScanOut1041;
wire [7:0] nOut16_18;
wire [7:0] nScanOut1042;
wire [7:0] nOut16_19;
wire [7:0] nScanOut1043;
wire [7:0] nOut16_20;
wire [7:0] nScanOut1044;
wire [7:0] nOut16_21;
wire [7:0] nScanOut1045;
wire [7:0] nOut16_22;
wire [7:0] nScanOut1046;
wire [7:0] nOut16_23;
wire [7:0] nScanOut1047;
wire [7:0] nOut16_24;
wire [7:0] nScanOut1048;
wire [7:0] nOut16_25;
wire [7:0] nScanOut1049;
wire [7:0] nOut16_26;
wire [7:0] nScanOut1050;
wire [7:0] nOut16_27;
wire [7:0] nScanOut1051;
wire [7:0] nOut16_28;
wire [7:0] nScanOut1052;
wire [7:0] nOut16_29;
wire [7:0] nScanOut1053;
wire [7:0] nOut16_30;
wire [7:0] nScanOut1054;
wire [7:0] nOut16_31;
wire [7:0] nScanOut1055;
wire [7:0] nOut16_32;
wire [7:0] nScanOut1056;
wire [7:0] nOut16_33;
wire [7:0] nScanOut1057;
wire [7:0] nOut16_34;
wire [7:0] nScanOut1058;
wire [7:0] nOut16_35;
wire [7:0] nScanOut1059;
wire [7:0] nOut16_36;
wire [7:0] nScanOut1060;
wire [7:0] nOut16_37;
wire [7:0] nScanOut1061;
wire [7:0] nOut16_38;
wire [7:0] nScanOut1062;
wire [7:0] nOut16_39;
wire [7:0] nScanOut1063;
wire [7:0] nOut16_40;
wire [7:0] nScanOut1064;
wire [7:0] nOut16_41;
wire [7:0] nScanOut1065;
wire [7:0] nOut16_42;
wire [7:0] nScanOut1066;
wire [7:0] nOut16_43;
wire [7:0] nScanOut1067;
wire [7:0] nOut16_44;
wire [7:0] nScanOut1068;
wire [7:0] nOut16_45;
wire [7:0] nScanOut1069;
wire [7:0] nOut16_46;
wire [7:0] nScanOut1070;
wire [7:0] nOut16_47;
wire [7:0] nScanOut1071;
wire [7:0] nOut16_48;
wire [7:0] nScanOut1072;
wire [7:0] nOut16_49;
wire [7:0] nScanOut1073;
wire [7:0] nOut16_50;
wire [7:0] nScanOut1074;
wire [7:0] nOut16_51;
wire [7:0] nScanOut1075;
wire [7:0] nOut16_52;
wire [7:0] nScanOut1076;
wire [7:0] nOut16_53;
wire [7:0] nScanOut1077;
wire [7:0] nOut16_54;
wire [7:0] nScanOut1078;
wire [7:0] nOut16_55;
wire [7:0] nScanOut1079;
wire [7:0] nOut16_56;
wire [7:0] nScanOut1080;
wire [7:0] nOut16_57;
wire [7:0] nScanOut1081;
wire [7:0] nOut16_58;
wire [7:0] nScanOut1082;
wire [7:0] nOut16_59;
wire [7:0] nScanOut1083;
wire [7:0] nOut16_60;
wire [7:0] nScanOut1084;
wire [7:0] nOut16_61;
wire [7:0] nScanOut1085;
wire [7:0] nOut16_62;
wire [7:0] nScanOut1086;
wire [7:0] nOut16_63;
wire [7:0] nScanOut1087;
wire [7:0] nOut17_0;
wire [7:0] nScanOut1088;
wire [7:0] nOut17_1;
wire [7:0] nScanOut1089;
wire [7:0] nOut17_2;
wire [7:0] nScanOut1090;
wire [7:0] nOut17_3;
wire [7:0] nScanOut1091;
wire [7:0] nOut17_4;
wire [7:0] nScanOut1092;
wire [7:0] nOut17_5;
wire [7:0] nScanOut1093;
wire [7:0] nOut17_6;
wire [7:0] nScanOut1094;
wire [7:0] nOut17_7;
wire [7:0] nScanOut1095;
wire [7:0] nOut17_8;
wire [7:0] nScanOut1096;
wire [7:0] nOut17_9;
wire [7:0] nScanOut1097;
wire [7:0] nOut17_10;
wire [7:0] nScanOut1098;
wire [7:0] nOut17_11;
wire [7:0] nScanOut1099;
wire [7:0] nOut17_12;
wire [7:0] nScanOut1100;
wire [7:0] nOut17_13;
wire [7:0] nScanOut1101;
wire [7:0] nOut17_14;
wire [7:0] nScanOut1102;
wire [7:0] nOut17_15;
wire [7:0] nScanOut1103;
wire [7:0] nOut17_16;
wire [7:0] nScanOut1104;
wire [7:0] nOut17_17;
wire [7:0] nScanOut1105;
wire [7:0] nOut17_18;
wire [7:0] nScanOut1106;
wire [7:0] nOut17_19;
wire [7:0] nScanOut1107;
wire [7:0] nOut17_20;
wire [7:0] nScanOut1108;
wire [7:0] nOut17_21;
wire [7:0] nScanOut1109;
wire [7:0] nOut17_22;
wire [7:0] nScanOut1110;
wire [7:0] nOut17_23;
wire [7:0] nScanOut1111;
wire [7:0] nOut17_24;
wire [7:0] nScanOut1112;
wire [7:0] nOut17_25;
wire [7:0] nScanOut1113;
wire [7:0] nOut17_26;
wire [7:0] nScanOut1114;
wire [7:0] nOut17_27;
wire [7:0] nScanOut1115;
wire [7:0] nOut17_28;
wire [7:0] nScanOut1116;
wire [7:0] nOut17_29;
wire [7:0] nScanOut1117;
wire [7:0] nOut17_30;
wire [7:0] nScanOut1118;
wire [7:0] nOut17_31;
wire [7:0] nScanOut1119;
wire [7:0] nOut17_32;
wire [7:0] nScanOut1120;
wire [7:0] nOut17_33;
wire [7:0] nScanOut1121;
wire [7:0] nOut17_34;
wire [7:0] nScanOut1122;
wire [7:0] nOut17_35;
wire [7:0] nScanOut1123;
wire [7:0] nOut17_36;
wire [7:0] nScanOut1124;
wire [7:0] nOut17_37;
wire [7:0] nScanOut1125;
wire [7:0] nOut17_38;
wire [7:0] nScanOut1126;
wire [7:0] nOut17_39;
wire [7:0] nScanOut1127;
wire [7:0] nOut17_40;
wire [7:0] nScanOut1128;
wire [7:0] nOut17_41;
wire [7:0] nScanOut1129;
wire [7:0] nOut17_42;
wire [7:0] nScanOut1130;
wire [7:0] nOut17_43;
wire [7:0] nScanOut1131;
wire [7:0] nOut17_44;
wire [7:0] nScanOut1132;
wire [7:0] nOut17_45;
wire [7:0] nScanOut1133;
wire [7:0] nOut17_46;
wire [7:0] nScanOut1134;
wire [7:0] nOut17_47;
wire [7:0] nScanOut1135;
wire [7:0] nOut17_48;
wire [7:0] nScanOut1136;
wire [7:0] nOut17_49;
wire [7:0] nScanOut1137;
wire [7:0] nOut17_50;
wire [7:0] nScanOut1138;
wire [7:0] nOut17_51;
wire [7:0] nScanOut1139;
wire [7:0] nOut17_52;
wire [7:0] nScanOut1140;
wire [7:0] nOut17_53;
wire [7:0] nScanOut1141;
wire [7:0] nOut17_54;
wire [7:0] nScanOut1142;
wire [7:0] nOut17_55;
wire [7:0] nScanOut1143;
wire [7:0] nOut17_56;
wire [7:0] nScanOut1144;
wire [7:0] nOut17_57;
wire [7:0] nScanOut1145;
wire [7:0] nOut17_58;
wire [7:0] nScanOut1146;
wire [7:0] nOut17_59;
wire [7:0] nScanOut1147;
wire [7:0] nOut17_60;
wire [7:0] nScanOut1148;
wire [7:0] nOut17_61;
wire [7:0] nScanOut1149;
wire [7:0] nOut17_62;
wire [7:0] nScanOut1150;
wire [7:0] nOut17_63;
wire [7:0] nScanOut1151;
wire [7:0] nOut18_0;
wire [7:0] nScanOut1152;
wire [7:0] nOut18_1;
wire [7:0] nScanOut1153;
wire [7:0] nOut18_2;
wire [7:0] nScanOut1154;
wire [7:0] nOut18_3;
wire [7:0] nScanOut1155;
wire [7:0] nOut18_4;
wire [7:0] nScanOut1156;
wire [7:0] nOut18_5;
wire [7:0] nScanOut1157;
wire [7:0] nOut18_6;
wire [7:0] nScanOut1158;
wire [7:0] nOut18_7;
wire [7:0] nScanOut1159;
wire [7:0] nOut18_8;
wire [7:0] nScanOut1160;
wire [7:0] nOut18_9;
wire [7:0] nScanOut1161;
wire [7:0] nOut18_10;
wire [7:0] nScanOut1162;
wire [7:0] nOut18_11;
wire [7:0] nScanOut1163;
wire [7:0] nOut18_12;
wire [7:0] nScanOut1164;
wire [7:0] nOut18_13;
wire [7:0] nScanOut1165;
wire [7:0] nOut18_14;
wire [7:0] nScanOut1166;
wire [7:0] nOut18_15;
wire [7:0] nScanOut1167;
wire [7:0] nOut18_16;
wire [7:0] nScanOut1168;
wire [7:0] nOut18_17;
wire [7:0] nScanOut1169;
wire [7:0] nOut18_18;
wire [7:0] nScanOut1170;
wire [7:0] nOut18_19;
wire [7:0] nScanOut1171;
wire [7:0] nOut18_20;
wire [7:0] nScanOut1172;
wire [7:0] nOut18_21;
wire [7:0] nScanOut1173;
wire [7:0] nOut18_22;
wire [7:0] nScanOut1174;
wire [7:0] nOut18_23;
wire [7:0] nScanOut1175;
wire [7:0] nOut18_24;
wire [7:0] nScanOut1176;
wire [7:0] nOut18_25;
wire [7:0] nScanOut1177;
wire [7:0] nOut18_26;
wire [7:0] nScanOut1178;
wire [7:0] nOut18_27;
wire [7:0] nScanOut1179;
wire [7:0] nOut18_28;
wire [7:0] nScanOut1180;
wire [7:0] nOut18_29;
wire [7:0] nScanOut1181;
wire [7:0] nOut18_30;
wire [7:0] nScanOut1182;
wire [7:0] nOut18_31;
wire [7:0] nScanOut1183;
wire [7:0] nOut18_32;
wire [7:0] nScanOut1184;
wire [7:0] nOut18_33;
wire [7:0] nScanOut1185;
wire [7:0] nOut18_34;
wire [7:0] nScanOut1186;
wire [7:0] nOut18_35;
wire [7:0] nScanOut1187;
wire [7:0] nOut18_36;
wire [7:0] nScanOut1188;
wire [7:0] nOut18_37;
wire [7:0] nScanOut1189;
wire [7:0] nOut18_38;
wire [7:0] nScanOut1190;
wire [7:0] nOut18_39;
wire [7:0] nScanOut1191;
wire [7:0] nOut18_40;
wire [7:0] nScanOut1192;
wire [7:0] nOut18_41;
wire [7:0] nScanOut1193;
wire [7:0] nOut18_42;
wire [7:0] nScanOut1194;
wire [7:0] nOut18_43;
wire [7:0] nScanOut1195;
wire [7:0] nOut18_44;
wire [7:0] nScanOut1196;
wire [7:0] nOut18_45;
wire [7:0] nScanOut1197;
wire [7:0] nOut18_46;
wire [7:0] nScanOut1198;
wire [7:0] nOut18_47;
wire [7:0] nScanOut1199;
wire [7:0] nOut18_48;
wire [7:0] nScanOut1200;
wire [7:0] nOut18_49;
wire [7:0] nScanOut1201;
wire [7:0] nOut18_50;
wire [7:0] nScanOut1202;
wire [7:0] nOut18_51;
wire [7:0] nScanOut1203;
wire [7:0] nOut18_52;
wire [7:0] nScanOut1204;
wire [7:0] nOut18_53;
wire [7:0] nScanOut1205;
wire [7:0] nOut18_54;
wire [7:0] nScanOut1206;
wire [7:0] nOut18_55;
wire [7:0] nScanOut1207;
wire [7:0] nOut18_56;
wire [7:0] nScanOut1208;
wire [7:0] nOut18_57;
wire [7:0] nScanOut1209;
wire [7:0] nOut18_58;
wire [7:0] nScanOut1210;
wire [7:0] nOut18_59;
wire [7:0] nScanOut1211;
wire [7:0] nOut18_60;
wire [7:0] nScanOut1212;
wire [7:0] nOut18_61;
wire [7:0] nScanOut1213;
wire [7:0] nOut18_62;
wire [7:0] nScanOut1214;
wire [7:0] nOut18_63;
wire [7:0] nScanOut1215;
wire [7:0] nOut19_0;
wire [7:0] nScanOut1216;
wire [7:0] nOut19_1;
wire [7:0] nScanOut1217;
wire [7:0] nOut19_2;
wire [7:0] nScanOut1218;
wire [7:0] nOut19_3;
wire [7:0] nScanOut1219;
wire [7:0] nOut19_4;
wire [7:0] nScanOut1220;
wire [7:0] nOut19_5;
wire [7:0] nScanOut1221;
wire [7:0] nOut19_6;
wire [7:0] nScanOut1222;
wire [7:0] nOut19_7;
wire [7:0] nScanOut1223;
wire [7:0] nOut19_8;
wire [7:0] nScanOut1224;
wire [7:0] nOut19_9;
wire [7:0] nScanOut1225;
wire [7:0] nOut19_10;
wire [7:0] nScanOut1226;
wire [7:0] nOut19_11;
wire [7:0] nScanOut1227;
wire [7:0] nOut19_12;
wire [7:0] nScanOut1228;
wire [7:0] nOut19_13;
wire [7:0] nScanOut1229;
wire [7:0] nOut19_14;
wire [7:0] nScanOut1230;
wire [7:0] nOut19_15;
wire [7:0] nScanOut1231;
wire [7:0] nOut19_16;
wire [7:0] nScanOut1232;
wire [7:0] nOut19_17;
wire [7:0] nScanOut1233;
wire [7:0] nOut19_18;
wire [7:0] nScanOut1234;
wire [7:0] nOut19_19;
wire [7:0] nScanOut1235;
wire [7:0] nOut19_20;
wire [7:0] nScanOut1236;
wire [7:0] nOut19_21;
wire [7:0] nScanOut1237;
wire [7:0] nOut19_22;
wire [7:0] nScanOut1238;
wire [7:0] nOut19_23;
wire [7:0] nScanOut1239;
wire [7:0] nOut19_24;
wire [7:0] nScanOut1240;
wire [7:0] nOut19_25;
wire [7:0] nScanOut1241;
wire [7:0] nOut19_26;
wire [7:0] nScanOut1242;
wire [7:0] nOut19_27;
wire [7:0] nScanOut1243;
wire [7:0] nOut19_28;
wire [7:0] nScanOut1244;
wire [7:0] nOut19_29;
wire [7:0] nScanOut1245;
wire [7:0] nOut19_30;
wire [7:0] nScanOut1246;
wire [7:0] nOut19_31;
wire [7:0] nScanOut1247;
wire [7:0] nOut19_32;
wire [7:0] nScanOut1248;
wire [7:0] nOut19_33;
wire [7:0] nScanOut1249;
wire [7:0] nOut19_34;
wire [7:0] nScanOut1250;
wire [7:0] nOut19_35;
wire [7:0] nScanOut1251;
wire [7:0] nOut19_36;
wire [7:0] nScanOut1252;
wire [7:0] nOut19_37;
wire [7:0] nScanOut1253;
wire [7:0] nOut19_38;
wire [7:0] nScanOut1254;
wire [7:0] nOut19_39;
wire [7:0] nScanOut1255;
wire [7:0] nOut19_40;
wire [7:0] nScanOut1256;
wire [7:0] nOut19_41;
wire [7:0] nScanOut1257;
wire [7:0] nOut19_42;
wire [7:0] nScanOut1258;
wire [7:0] nOut19_43;
wire [7:0] nScanOut1259;
wire [7:0] nOut19_44;
wire [7:0] nScanOut1260;
wire [7:0] nOut19_45;
wire [7:0] nScanOut1261;
wire [7:0] nOut19_46;
wire [7:0] nScanOut1262;
wire [7:0] nOut19_47;
wire [7:0] nScanOut1263;
wire [7:0] nOut19_48;
wire [7:0] nScanOut1264;
wire [7:0] nOut19_49;
wire [7:0] nScanOut1265;
wire [7:0] nOut19_50;
wire [7:0] nScanOut1266;
wire [7:0] nOut19_51;
wire [7:0] nScanOut1267;
wire [7:0] nOut19_52;
wire [7:0] nScanOut1268;
wire [7:0] nOut19_53;
wire [7:0] nScanOut1269;
wire [7:0] nOut19_54;
wire [7:0] nScanOut1270;
wire [7:0] nOut19_55;
wire [7:0] nScanOut1271;
wire [7:0] nOut19_56;
wire [7:0] nScanOut1272;
wire [7:0] nOut19_57;
wire [7:0] nScanOut1273;
wire [7:0] nOut19_58;
wire [7:0] nScanOut1274;
wire [7:0] nOut19_59;
wire [7:0] nScanOut1275;
wire [7:0] nOut19_60;
wire [7:0] nScanOut1276;
wire [7:0] nOut19_61;
wire [7:0] nScanOut1277;
wire [7:0] nOut19_62;
wire [7:0] nScanOut1278;
wire [7:0] nOut19_63;
wire [7:0] nScanOut1279;
wire [7:0] nOut20_0;
wire [7:0] nScanOut1280;
wire [7:0] nOut20_1;
wire [7:0] nScanOut1281;
wire [7:0] nOut20_2;
wire [7:0] nScanOut1282;
wire [7:0] nOut20_3;
wire [7:0] nScanOut1283;
wire [7:0] nOut20_4;
wire [7:0] nScanOut1284;
wire [7:0] nOut20_5;
wire [7:0] nScanOut1285;
wire [7:0] nOut20_6;
wire [7:0] nScanOut1286;
wire [7:0] nOut20_7;
wire [7:0] nScanOut1287;
wire [7:0] nOut20_8;
wire [7:0] nScanOut1288;
wire [7:0] nOut20_9;
wire [7:0] nScanOut1289;
wire [7:0] nOut20_10;
wire [7:0] nScanOut1290;
wire [7:0] nOut20_11;
wire [7:0] nScanOut1291;
wire [7:0] nOut20_12;
wire [7:0] nScanOut1292;
wire [7:0] nOut20_13;
wire [7:0] nScanOut1293;
wire [7:0] nOut20_14;
wire [7:0] nScanOut1294;
wire [7:0] nOut20_15;
wire [7:0] nScanOut1295;
wire [7:0] nOut20_16;
wire [7:0] nScanOut1296;
wire [7:0] nOut20_17;
wire [7:0] nScanOut1297;
wire [7:0] nOut20_18;
wire [7:0] nScanOut1298;
wire [7:0] nOut20_19;
wire [7:0] nScanOut1299;
wire [7:0] nOut20_20;
wire [7:0] nScanOut1300;
wire [7:0] nOut20_21;
wire [7:0] nScanOut1301;
wire [7:0] nOut20_22;
wire [7:0] nScanOut1302;
wire [7:0] nOut20_23;
wire [7:0] nScanOut1303;
wire [7:0] nOut20_24;
wire [7:0] nScanOut1304;
wire [7:0] nOut20_25;
wire [7:0] nScanOut1305;
wire [7:0] nOut20_26;
wire [7:0] nScanOut1306;
wire [7:0] nOut20_27;
wire [7:0] nScanOut1307;
wire [7:0] nOut20_28;
wire [7:0] nScanOut1308;
wire [7:0] nOut20_29;
wire [7:0] nScanOut1309;
wire [7:0] nOut20_30;
wire [7:0] nScanOut1310;
wire [7:0] nOut20_31;
wire [7:0] nScanOut1311;
wire [7:0] nOut20_32;
wire [7:0] nScanOut1312;
wire [7:0] nOut20_33;
wire [7:0] nScanOut1313;
wire [7:0] nOut20_34;
wire [7:0] nScanOut1314;
wire [7:0] nOut20_35;
wire [7:0] nScanOut1315;
wire [7:0] nOut20_36;
wire [7:0] nScanOut1316;
wire [7:0] nOut20_37;
wire [7:0] nScanOut1317;
wire [7:0] nOut20_38;
wire [7:0] nScanOut1318;
wire [7:0] nOut20_39;
wire [7:0] nScanOut1319;
wire [7:0] nOut20_40;
wire [7:0] nScanOut1320;
wire [7:0] nOut20_41;
wire [7:0] nScanOut1321;
wire [7:0] nOut20_42;
wire [7:0] nScanOut1322;
wire [7:0] nOut20_43;
wire [7:0] nScanOut1323;
wire [7:0] nOut20_44;
wire [7:0] nScanOut1324;
wire [7:0] nOut20_45;
wire [7:0] nScanOut1325;
wire [7:0] nOut20_46;
wire [7:0] nScanOut1326;
wire [7:0] nOut20_47;
wire [7:0] nScanOut1327;
wire [7:0] nOut20_48;
wire [7:0] nScanOut1328;
wire [7:0] nOut20_49;
wire [7:0] nScanOut1329;
wire [7:0] nOut20_50;
wire [7:0] nScanOut1330;
wire [7:0] nOut20_51;
wire [7:0] nScanOut1331;
wire [7:0] nOut20_52;
wire [7:0] nScanOut1332;
wire [7:0] nOut20_53;
wire [7:0] nScanOut1333;
wire [7:0] nOut20_54;
wire [7:0] nScanOut1334;
wire [7:0] nOut20_55;
wire [7:0] nScanOut1335;
wire [7:0] nOut20_56;
wire [7:0] nScanOut1336;
wire [7:0] nOut20_57;
wire [7:0] nScanOut1337;
wire [7:0] nOut20_58;
wire [7:0] nScanOut1338;
wire [7:0] nOut20_59;
wire [7:0] nScanOut1339;
wire [7:0] nOut20_60;
wire [7:0] nScanOut1340;
wire [7:0] nOut20_61;
wire [7:0] nScanOut1341;
wire [7:0] nOut20_62;
wire [7:0] nScanOut1342;
wire [7:0] nOut20_63;
wire [7:0] nScanOut1343;
wire [7:0] nOut21_0;
wire [7:0] nScanOut1344;
wire [7:0] nOut21_1;
wire [7:0] nScanOut1345;
wire [7:0] nOut21_2;
wire [7:0] nScanOut1346;
wire [7:0] nOut21_3;
wire [7:0] nScanOut1347;
wire [7:0] nOut21_4;
wire [7:0] nScanOut1348;
wire [7:0] nOut21_5;
wire [7:0] nScanOut1349;
wire [7:0] nOut21_6;
wire [7:0] nScanOut1350;
wire [7:0] nOut21_7;
wire [7:0] nScanOut1351;
wire [7:0] nOut21_8;
wire [7:0] nScanOut1352;
wire [7:0] nOut21_9;
wire [7:0] nScanOut1353;
wire [7:0] nOut21_10;
wire [7:0] nScanOut1354;
wire [7:0] nOut21_11;
wire [7:0] nScanOut1355;
wire [7:0] nOut21_12;
wire [7:0] nScanOut1356;
wire [7:0] nOut21_13;
wire [7:0] nScanOut1357;
wire [7:0] nOut21_14;
wire [7:0] nScanOut1358;
wire [7:0] nOut21_15;
wire [7:0] nScanOut1359;
wire [7:0] nOut21_16;
wire [7:0] nScanOut1360;
wire [7:0] nOut21_17;
wire [7:0] nScanOut1361;
wire [7:0] nOut21_18;
wire [7:0] nScanOut1362;
wire [7:0] nOut21_19;
wire [7:0] nScanOut1363;
wire [7:0] nOut21_20;
wire [7:0] nScanOut1364;
wire [7:0] nOut21_21;
wire [7:0] nScanOut1365;
wire [7:0] nOut21_22;
wire [7:0] nScanOut1366;
wire [7:0] nOut21_23;
wire [7:0] nScanOut1367;
wire [7:0] nOut21_24;
wire [7:0] nScanOut1368;
wire [7:0] nOut21_25;
wire [7:0] nScanOut1369;
wire [7:0] nOut21_26;
wire [7:0] nScanOut1370;
wire [7:0] nOut21_27;
wire [7:0] nScanOut1371;
wire [7:0] nOut21_28;
wire [7:0] nScanOut1372;
wire [7:0] nOut21_29;
wire [7:0] nScanOut1373;
wire [7:0] nOut21_30;
wire [7:0] nScanOut1374;
wire [7:0] nOut21_31;
wire [7:0] nScanOut1375;
wire [7:0] nOut21_32;
wire [7:0] nScanOut1376;
wire [7:0] nOut21_33;
wire [7:0] nScanOut1377;
wire [7:0] nOut21_34;
wire [7:0] nScanOut1378;
wire [7:0] nOut21_35;
wire [7:0] nScanOut1379;
wire [7:0] nOut21_36;
wire [7:0] nScanOut1380;
wire [7:0] nOut21_37;
wire [7:0] nScanOut1381;
wire [7:0] nOut21_38;
wire [7:0] nScanOut1382;
wire [7:0] nOut21_39;
wire [7:0] nScanOut1383;
wire [7:0] nOut21_40;
wire [7:0] nScanOut1384;
wire [7:0] nOut21_41;
wire [7:0] nScanOut1385;
wire [7:0] nOut21_42;
wire [7:0] nScanOut1386;
wire [7:0] nOut21_43;
wire [7:0] nScanOut1387;
wire [7:0] nOut21_44;
wire [7:0] nScanOut1388;
wire [7:0] nOut21_45;
wire [7:0] nScanOut1389;
wire [7:0] nOut21_46;
wire [7:0] nScanOut1390;
wire [7:0] nOut21_47;
wire [7:0] nScanOut1391;
wire [7:0] nOut21_48;
wire [7:0] nScanOut1392;
wire [7:0] nOut21_49;
wire [7:0] nScanOut1393;
wire [7:0] nOut21_50;
wire [7:0] nScanOut1394;
wire [7:0] nOut21_51;
wire [7:0] nScanOut1395;
wire [7:0] nOut21_52;
wire [7:0] nScanOut1396;
wire [7:0] nOut21_53;
wire [7:0] nScanOut1397;
wire [7:0] nOut21_54;
wire [7:0] nScanOut1398;
wire [7:0] nOut21_55;
wire [7:0] nScanOut1399;
wire [7:0] nOut21_56;
wire [7:0] nScanOut1400;
wire [7:0] nOut21_57;
wire [7:0] nScanOut1401;
wire [7:0] nOut21_58;
wire [7:0] nScanOut1402;
wire [7:0] nOut21_59;
wire [7:0] nScanOut1403;
wire [7:0] nOut21_60;
wire [7:0] nScanOut1404;
wire [7:0] nOut21_61;
wire [7:0] nScanOut1405;
wire [7:0] nOut21_62;
wire [7:0] nScanOut1406;
wire [7:0] nOut21_63;
wire [7:0] nScanOut1407;
wire [7:0] nOut22_0;
wire [7:0] nScanOut1408;
wire [7:0] nOut22_1;
wire [7:0] nScanOut1409;
wire [7:0] nOut22_2;
wire [7:0] nScanOut1410;
wire [7:0] nOut22_3;
wire [7:0] nScanOut1411;
wire [7:0] nOut22_4;
wire [7:0] nScanOut1412;
wire [7:0] nOut22_5;
wire [7:0] nScanOut1413;
wire [7:0] nOut22_6;
wire [7:0] nScanOut1414;
wire [7:0] nOut22_7;
wire [7:0] nScanOut1415;
wire [7:0] nOut22_8;
wire [7:0] nScanOut1416;
wire [7:0] nOut22_9;
wire [7:0] nScanOut1417;
wire [7:0] nOut22_10;
wire [7:0] nScanOut1418;
wire [7:0] nOut22_11;
wire [7:0] nScanOut1419;
wire [7:0] nOut22_12;
wire [7:0] nScanOut1420;
wire [7:0] nOut22_13;
wire [7:0] nScanOut1421;
wire [7:0] nOut22_14;
wire [7:0] nScanOut1422;
wire [7:0] nOut22_15;
wire [7:0] nScanOut1423;
wire [7:0] nOut22_16;
wire [7:0] nScanOut1424;
wire [7:0] nOut22_17;
wire [7:0] nScanOut1425;
wire [7:0] nOut22_18;
wire [7:0] nScanOut1426;
wire [7:0] nOut22_19;
wire [7:0] nScanOut1427;
wire [7:0] nOut22_20;
wire [7:0] nScanOut1428;
wire [7:0] nOut22_21;
wire [7:0] nScanOut1429;
wire [7:0] nOut22_22;
wire [7:0] nScanOut1430;
wire [7:0] nOut22_23;
wire [7:0] nScanOut1431;
wire [7:0] nOut22_24;
wire [7:0] nScanOut1432;
wire [7:0] nOut22_25;
wire [7:0] nScanOut1433;
wire [7:0] nOut22_26;
wire [7:0] nScanOut1434;
wire [7:0] nOut22_27;
wire [7:0] nScanOut1435;
wire [7:0] nOut22_28;
wire [7:0] nScanOut1436;
wire [7:0] nOut22_29;
wire [7:0] nScanOut1437;
wire [7:0] nOut22_30;
wire [7:0] nScanOut1438;
wire [7:0] nOut22_31;
wire [7:0] nScanOut1439;
wire [7:0] nOut22_32;
wire [7:0] nScanOut1440;
wire [7:0] nOut22_33;
wire [7:0] nScanOut1441;
wire [7:0] nOut22_34;
wire [7:0] nScanOut1442;
wire [7:0] nOut22_35;
wire [7:0] nScanOut1443;
wire [7:0] nOut22_36;
wire [7:0] nScanOut1444;
wire [7:0] nOut22_37;
wire [7:0] nScanOut1445;
wire [7:0] nOut22_38;
wire [7:0] nScanOut1446;
wire [7:0] nOut22_39;
wire [7:0] nScanOut1447;
wire [7:0] nOut22_40;
wire [7:0] nScanOut1448;
wire [7:0] nOut22_41;
wire [7:0] nScanOut1449;
wire [7:0] nOut22_42;
wire [7:0] nScanOut1450;
wire [7:0] nOut22_43;
wire [7:0] nScanOut1451;
wire [7:0] nOut22_44;
wire [7:0] nScanOut1452;
wire [7:0] nOut22_45;
wire [7:0] nScanOut1453;
wire [7:0] nOut22_46;
wire [7:0] nScanOut1454;
wire [7:0] nOut22_47;
wire [7:0] nScanOut1455;
wire [7:0] nOut22_48;
wire [7:0] nScanOut1456;
wire [7:0] nOut22_49;
wire [7:0] nScanOut1457;
wire [7:0] nOut22_50;
wire [7:0] nScanOut1458;
wire [7:0] nOut22_51;
wire [7:0] nScanOut1459;
wire [7:0] nOut22_52;
wire [7:0] nScanOut1460;
wire [7:0] nOut22_53;
wire [7:0] nScanOut1461;
wire [7:0] nOut22_54;
wire [7:0] nScanOut1462;
wire [7:0] nOut22_55;
wire [7:0] nScanOut1463;
wire [7:0] nOut22_56;
wire [7:0] nScanOut1464;
wire [7:0] nOut22_57;
wire [7:0] nScanOut1465;
wire [7:0] nOut22_58;
wire [7:0] nScanOut1466;
wire [7:0] nOut22_59;
wire [7:0] nScanOut1467;
wire [7:0] nOut22_60;
wire [7:0] nScanOut1468;
wire [7:0] nOut22_61;
wire [7:0] nScanOut1469;
wire [7:0] nOut22_62;
wire [7:0] nScanOut1470;
wire [7:0] nOut22_63;
wire [7:0] nScanOut1471;
wire [7:0] nOut23_0;
wire [7:0] nScanOut1472;
wire [7:0] nOut23_1;
wire [7:0] nScanOut1473;
wire [7:0] nOut23_2;
wire [7:0] nScanOut1474;
wire [7:0] nOut23_3;
wire [7:0] nScanOut1475;
wire [7:0] nOut23_4;
wire [7:0] nScanOut1476;
wire [7:0] nOut23_5;
wire [7:0] nScanOut1477;
wire [7:0] nOut23_6;
wire [7:0] nScanOut1478;
wire [7:0] nOut23_7;
wire [7:0] nScanOut1479;
wire [7:0] nOut23_8;
wire [7:0] nScanOut1480;
wire [7:0] nOut23_9;
wire [7:0] nScanOut1481;
wire [7:0] nOut23_10;
wire [7:0] nScanOut1482;
wire [7:0] nOut23_11;
wire [7:0] nScanOut1483;
wire [7:0] nOut23_12;
wire [7:0] nScanOut1484;
wire [7:0] nOut23_13;
wire [7:0] nScanOut1485;
wire [7:0] nOut23_14;
wire [7:0] nScanOut1486;
wire [7:0] nOut23_15;
wire [7:0] nScanOut1487;
wire [7:0] nOut23_16;
wire [7:0] nScanOut1488;
wire [7:0] nOut23_17;
wire [7:0] nScanOut1489;
wire [7:0] nOut23_18;
wire [7:0] nScanOut1490;
wire [7:0] nOut23_19;
wire [7:0] nScanOut1491;
wire [7:0] nOut23_20;
wire [7:0] nScanOut1492;
wire [7:0] nOut23_21;
wire [7:0] nScanOut1493;
wire [7:0] nOut23_22;
wire [7:0] nScanOut1494;
wire [7:0] nOut23_23;
wire [7:0] nScanOut1495;
wire [7:0] nOut23_24;
wire [7:0] nScanOut1496;
wire [7:0] nOut23_25;
wire [7:0] nScanOut1497;
wire [7:0] nOut23_26;
wire [7:0] nScanOut1498;
wire [7:0] nOut23_27;
wire [7:0] nScanOut1499;
wire [7:0] nOut23_28;
wire [7:0] nScanOut1500;
wire [7:0] nOut23_29;
wire [7:0] nScanOut1501;
wire [7:0] nOut23_30;
wire [7:0] nScanOut1502;
wire [7:0] nOut23_31;
wire [7:0] nScanOut1503;
wire [7:0] nOut23_32;
wire [7:0] nScanOut1504;
wire [7:0] nOut23_33;
wire [7:0] nScanOut1505;
wire [7:0] nOut23_34;
wire [7:0] nScanOut1506;
wire [7:0] nOut23_35;
wire [7:0] nScanOut1507;
wire [7:0] nOut23_36;
wire [7:0] nScanOut1508;
wire [7:0] nOut23_37;
wire [7:0] nScanOut1509;
wire [7:0] nOut23_38;
wire [7:0] nScanOut1510;
wire [7:0] nOut23_39;
wire [7:0] nScanOut1511;
wire [7:0] nOut23_40;
wire [7:0] nScanOut1512;
wire [7:0] nOut23_41;
wire [7:0] nScanOut1513;
wire [7:0] nOut23_42;
wire [7:0] nScanOut1514;
wire [7:0] nOut23_43;
wire [7:0] nScanOut1515;
wire [7:0] nOut23_44;
wire [7:0] nScanOut1516;
wire [7:0] nOut23_45;
wire [7:0] nScanOut1517;
wire [7:0] nOut23_46;
wire [7:0] nScanOut1518;
wire [7:0] nOut23_47;
wire [7:0] nScanOut1519;
wire [7:0] nOut23_48;
wire [7:0] nScanOut1520;
wire [7:0] nOut23_49;
wire [7:0] nScanOut1521;
wire [7:0] nOut23_50;
wire [7:0] nScanOut1522;
wire [7:0] nOut23_51;
wire [7:0] nScanOut1523;
wire [7:0] nOut23_52;
wire [7:0] nScanOut1524;
wire [7:0] nOut23_53;
wire [7:0] nScanOut1525;
wire [7:0] nOut23_54;
wire [7:0] nScanOut1526;
wire [7:0] nOut23_55;
wire [7:0] nScanOut1527;
wire [7:0] nOut23_56;
wire [7:0] nScanOut1528;
wire [7:0] nOut23_57;
wire [7:0] nScanOut1529;
wire [7:0] nOut23_58;
wire [7:0] nScanOut1530;
wire [7:0] nOut23_59;
wire [7:0] nScanOut1531;
wire [7:0] nOut23_60;
wire [7:0] nScanOut1532;
wire [7:0] nOut23_61;
wire [7:0] nScanOut1533;
wire [7:0] nOut23_62;
wire [7:0] nScanOut1534;
wire [7:0] nOut23_63;
wire [7:0] nScanOut1535;
wire [7:0] nOut24_0;
wire [7:0] nScanOut1536;
wire [7:0] nOut24_1;
wire [7:0] nScanOut1537;
wire [7:0] nOut24_2;
wire [7:0] nScanOut1538;
wire [7:0] nOut24_3;
wire [7:0] nScanOut1539;
wire [7:0] nOut24_4;
wire [7:0] nScanOut1540;
wire [7:0] nOut24_5;
wire [7:0] nScanOut1541;
wire [7:0] nOut24_6;
wire [7:0] nScanOut1542;
wire [7:0] nOut24_7;
wire [7:0] nScanOut1543;
wire [7:0] nOut24_8;
wire [7:0] nScanOut1544;
wire [7:0] nOut24_9;
wire [7:0] nScanOut1545;
wire [7:0] nOut24_10;
wire [7:0] nScanOut1546;
wire [7:0] nOut24_11;
wire [7:0] nScanOut1547;
wire [7:0] nOut24_12;
wire [7:0] nScanOut1548;
wire [7:0] nOut24_13;
wire [7:0] nScanOut1549;
wire [7:0] nOut24_14;
wire [7:0] nScanOut1550;
wire [7:0] nOut24_15;
wire [7:0] nScanOut1551;
wire [7:0] nOut24_16;
wire [7:0] nScanOut1552;
wire [7:0] nOut24_17;
wire [7:0] nScanOut1553;
wire [7:0] nOut24_18;
wire [7:0] nScanOut1554;
wire [7:0] nOut24_19;
wire [7:0] nScanOut1555;
wire [7:0] nOut24_20;
wire [7:0] nScanOut1556;
wire [7:0] nOut24_21;
wire [7:0] nScanOut1557;
wire [7:0] nOut24_22;
wire [7:0] nScanOut1558;
wire [7:0] nOut24_23;
wire [7:0] nScanOut1559;
wire [7:0] nOut24_24;
wire [7:0] nScanOut1560;
wire [7:0] nOut24_25;
wire [7:0] nScanOut1561;
wire [7:0] nOut24_26;
wire [7:0] nScanOut1562;
wire [7:0] nOut24_27;
wire [7:0] nScanOut1563;
wire [7:0] nOut24_28;
wire [7:0] nScanOut1564;
wire [7:0] nOut24_29;
wire [7:0] nScanOut1565;
wire [7:0] nOut24_30;
wire [7:0] nScanOut1566;
wire [7:0] nOut24_31;
wire [7:0] nScanOut1567;
wire [7:0] nOut24_32;
wire [7:0] nScanOut1568;
wire [7:0] nOut24_33;
wire [7:0] nScanOut1569;
wire [7:0] nOut24_34;
wire [7:0] nScanOut1570;
wire [7:0] nOut24_35;
wire [7:0] nScanOut1571;
wire [7:0] nOut24_36;
wire [7:0] nScanOut1572;
wire [7:0] nOut24_37;
wire [7:0] nScanOut1573;
wire [7:0] nOut24_38;
wire [7:0] nScanOut1574;
wire [7:0] nOut24_39;
wire [7:0] nScanOut1575;
wire [7:0] nOut24_40;
wire [7:0] nScanOut1576;
wire [7:0] nOut24_41;
wire [7:0] nScanOut1577;
wire [7:0] nOut24_42;
wire [7:0] nScanOut1578;
wire [7:0] nOut24_43;
wire [7:0] nScanOut1579;
wire [7:0] nOut24_44;
wire [7:0] nScanOut1580;
wire [7:0] nOut24_45;
wire [7:0] nScanOut1581;
wire [7:0] nOut24_46;
wire [7:0] nScanOut1582;
wire [7:0] nOut24_47;
wire [7:0] nScanOut1583;
wire [7:0] nOut24_48;
wire [7:0] nScanOut1584;
wire [7:0] nOut24_49;
wire [7:0] nScanOut1585;
wire [7:0] nOut24_50;
wire [7:0] nScanOut1586;
wire [7:0] nOut24_51;
wire [7:0] nScanOut1587;
wire [7:0] nOut24_52;
wire [7:0] nScanOut1588;
wire [7:0] nOut24_53;
wire [7:0] nScanOut1589;
wire [7:0] nOut24_54;
wire [7:0] nScanOut1590;
wire [7:0] nOut24_55;
wire [7:0] nScanOut1591;
wire [7:0] nOut24_56;
wire [7:0] nScanOut1592;
wire [7:0] nOut24_57;
wire [7:0] nScanOut1593;
wire [7:0] nOut24_58;
wire [7:0] nScanOut1594;
wire [7:0] nOut24_59;
wire [7:0] nScanOut1595;
wire [7:0] nOut24_60;
wire [7:0] nScanOut1596;
wire [7:0] nOut24_61;
wire [7:0] nScanOut1597;
wire [7:0] nOut24_62;
wire [7:0] nScanOut1598;
wire [7:0] nOut24_63;
wire [7:0] nScanOut1599;
wire [7:0] nOut25_0;
wire [7:0] nScanOut1600;
wire [7:0] nOut25_1;
wire [7:0] nScanOut1601;
wire [7:0] nOut25_2;
wire [7:0] nScanOut1602;
wire [7:0] nOut25_3;
wire [7:0] nScanOut1603;
wire [7:0] nOut25_4;
wire [7:0] nScanOut1604;
wire [7:0] nOut25_5;
wire [7:0] nScanOut1605;
wire [7:0] nOut25_6;
wire [7:0] nScanOut1606;
wire [7:0] nOut25_7;
wire [7:0] nScanOut1607;
wire [7:0] nOut25_8;
wire [7:0] nScanOut1608;
wire [7:0] nOut25_9;
wire [7:0] nScanOut1609;
wire [7:0] nOut25_10;
wire [7:0] nScanOut1610;
wire [7:0] nOut25_11;
wire [7:0] nScanOut1611;
wire [7:0] nOut25_12;
wire [7:0] nScanOut1612;
wire [7:0] nOut25_13;
wire [7:0] nScanOut1613;
wire [7:0] nOut25_14;
wire [7:0] nScanOut1614;
wire [7:0] nOut25_15;
wire [7:0] nScanOut1615;
wire [7:0] nOut25_16;
wire [7:0] nScanOut1616;
wire [7:0] nOut25_17;
wire [7:0] nScanOut1617;
wire [7:0] nOut25_18;
wire [7:0] nScanOut1618;
wire [7:0] nOut25_19;
wire [7:0] nScanOut1619;
wire [7:0] nOut25_20;
wire [7:0] nScanOut1620;
wire [7:0] nOut25_21;
wire [7:0] nScanOut1621;
wire [7:0] nOut25_22;
wire [7:0] nScanOut1622;
wire [7:0] nOut25_23;
wire [7:0] nScanOut1623;
wire [7:0] nOut25_24;
wire [7:0] nScanOut1624;
wire [7:0] nOut25_25;
wire [7:0] nScanOut1625;
wire [7:0] nOut25_26;
wire [7:0] nScanOut1626;
wire [7:0] nOut25_27;
wire [7:0] nScanOut1627;
wire [7:0] nOut25_28;
wire [7:0] nScanOut1628;
wire [7:0] nOut25_29;
wire [7:0] nScanOut1629;
wire [7:0] nOut25_30;
wire [7:0] nScanOut1630;
wire [7:0] nOut25_31;
wire [7:0] nScanOut1631;
wire [7:0] nOut25_32;
wire [7:0] nScanOut1632;
wire [7:0] nOut25_33;
wire [7:0] nScanOut1633;
wire [7:0] nOut25_34;
wire [7:0] nScanOut1634;
wire [7:0] nOut25_35;
wire [7:0] nScanOut1635;
wire [7:0] nOut25_36;
wire [7:0] nScanOut1636;
wire [7:0] nOut25_37;
wire [7:0] nScanOut1637;
wire [7:0] nOut25_38;
wire [7:0] nScanOut1638;
wire [7:0] nOut25_39;
wire [7:0] nScanOut1639;
wire [7:0] nOut25_40;
wire [7:0] nScanOut1640;
wire [7:0] nOut25_41;
wire [7:0] nScanOut1641;
wire [7:0] nOut25_42;
wire [7:0] nScanOut1642;
wire [7:0] nOut25_43;
wire [7:0] nScanOut1643;
wire [7:0] nOut25_44;
wire [7:0] nScanOut1644;
wire [7:0] nOut25_45;
wire [7:0] nScanOut1645;
wire [7:0] nOut25_46;
wire [7:0] nScanOut1646;
wire [7:0] nOut25_47;
wire [7:0] nScanOut1647;
wire [7:0] nOut25_48;
wire [7:0] nScanOut1648;
wire [7:0] nOut25_49;
wire [7:0] nScanOut1649;
wire [7:0] nOut25_50;
wire [7:0] nScanOut1650;
wire [7:0] nOut25_51;
wire [7:0] nScanOut1651;
wire [7:0] nOut25_52;
wire [7:0] nScanOut1652;
wire [7:0] nOut25_53;
wire [7:0] nScanOut1653;
wire [7:0] nOut25_54;
wire [7:0] nScanOut1654;
wire [7:0] nOut25_55;
wire [7:0] nScanOut1655;
wire [7:0] nOut25_56;
wire [7:0] nScanOut1656;
wire [7:0] nOut25_57;
wire [7:0] nScanOut1657;
wire [7:0] nOut25_58;
wire [7:0] nScanOut1658;
wire [7:0] nOut25_59;
wire [7:0] nScanOut1659;
wire [7:0] nOut25_60;
wire [7:0] nScanOut1660;
wire [7:0] nOut25_61;
wire [7:0] nScanOut1661;
wire [7:0] nOut25_62;
wire [7:0] nScanOut1662;
wire [7:0] nOut25_63;
wire [7:0] nScanOut1663;
wire [7:0] nOut26_0;
wire [7:0] nScanOut1664;
wire [7:0] nOut26_1;
wire [7:0] nScanOut1665;
wire [7:0] nOut26_2;
wire [7:0] nScanOut1666;
wire [7:0] nOut26_3;
wire [7:0] nScanOut1667;
wire [7:0] nOut26_4;
wire [7:0] nScanOut1668;
wire [7:0] nOut26_5;
wire [7:0] nScanOut1669;
wire [7:0] nOut26_6;
wire [7:0] nScanOut1670;
wire [7:0] nOut26_7;
wire [7:0] nScanOut1671;
wire [7:0] nOut26_8;
wire [7:0] nScanOut1672;
wire [7:0] nOut26_9;
wire [7:0] nScanOut1673;
wire [7:0] nOut26_10;
wire [7:0] nScanOut1674;
wire [7:0] nOut26_11;
wire [7:0] nScanOut1675;
wire [7:0] nOut26_12;
wire [7:0] nScanOut1676;
wire [7:0] nOut26_13;
wire [7:0] nScanOut1677;
wire [7:0] nOut26_14;
wire [7:0] nScanOut1678;
wire [7:0] nOut26_15;
wire [7:0] nScanOut1679;
wire [7:0] nOut26_16;
wire [7:0] nScanOut1680;
wire [7:0] nOut26_17;
wire [7:0] nScanOut1681;
wire [7:0] nOut26_18;
wire [7:0] nScanOut1682;
wire [7:0] nOut26_19;
wire [7:0] nScanOut1683;
wire [7:0] nOut26_20;
wire [7:0] nScanOut1684;
wire [7:0] nOut26_21;
wire [7:0] nScanOut1685;
wire [7:0] nOut26_22;
wire [7:0] nScanOut1686;
wire [7:0] nOut26_23;
wire [7:0] nScanOut1687;
wire [7:0] nOut26_24;
wire [7:0] nScanOut1688;
wire [7:0] nOut26_25;
wire [7:0] nScanOut1689;
wire [7:0] nOut26_26;
wire [7:0] nScanOut1690;
wire [7:0] nOut26_27;
wire [7:0] nScanOut1691;
wire [7:0] nOut26_28;
wire [7:0] nScanOut1692;
wire [7:0] nOut26_29;
wire [7:0] nScanOut1693;
wire [7:0] nOut26_30;
wire [7:0] nScanOut1694;
wire [7:0] nOut26_31;
wire [7:0] nScanOut1695;
wire [7:0] nOut26_32;
wire [7:0] nScanOut1696;
wire [7:0] nOut26_33;
wire [7:0] nScanOut1697;
wire [7:0] nOut26_34;
wire [7:0] nScanOut1698;
wire [7:0] nOut26_35;
wire [7:0] nScanOut1699;
wire [7:0] nOut26_36;
wire [7:0] nScanOut1700;
wire [7:0] nOut26_37;
wire [7:0] nScanOut1701;
wire [7:0] nOut26_38;
wire [7:0] nScanOut1702;
wire [7:0] nOut26_39;
wire [7:0] nScanOut1703;
wire [7:0] nOut26_40;
wire [7:0] nScanOut1704;
wire [7:0] nOut26_41;
wire [7:0] nScanOut1705;
wire [7:0] nOut26_42;
wire [7:0] nScanOut1706;
wire [7:0] nOut26_43;
wire [7:0] nScanOut1707;
wire [7:0] nOut26_44;
wire [7:0] nScanOut1708;
wire [7:0] nOut26_45;
wire [7:0] nScanOut1709;
wire [7:0] nOut26_46;
wire [7:0] nScanOut1710;
wire [7:0] nOut26_47;
wire [7:0] nScanOut1711;
wire [7:0] nOut26_48;
wire [7:0] nScanOut1712;
wire [7:0] nOut26_49;
wire [7:0] nScanOut1713;
wire [7:0] nOut26_50;
wire [7:0] nScanOut1714;
wire [7:0] nOut26_51;
wire [7:0] nScanOut1715;
wire [7:0] nOut26_52;
wire [7:0] nScanOut1716;
wire [7:0] nOut26_53;
wire [7:0] nScanOut1717;
wire [7:0] nOut26_54;
wire [7:0] nScanOut1718;
wire [7:0] nOut26_55;
wire [7:0] nScanOut1719;
wire [7:0] nOut26_56;
wire [7:0] nScanOut1720;
wire [7:0] nOut26_57;
wire [7:0] nScanOut1721;
wire [7:0] nOut26_58;
wire [7:0] nScanOut1722;
wire [7:0] nOut26_59;
wire [7:0] nScanOut1723;
wire [7:0] nOut26_60;
wire [7:0] nScanOut1724;
wire [7:0] nOut26_61;
wire [7:0] nScanOut1725;
wire [7:0] nOut26_62;
wire [7:0] nScanOut1726;
wire [7:0] nOut26_63;
wire [7:0] nScanOut1727;
wire [7:0] nOut27_0;
wire [7:0] nScanOut1728;
wire [7:0] nOut27_1;
wire [7:0] nScanOut1729;
wire [7:0] nOut27_2;
wire [7:0] nScanOut1730;
wire [7:0] nOut27_3;
wire [7:0] nScanOut1731;
wire [7:0] nOut27_4;
wire [7:0] nScanOut1732;
wire [7:0] nOut27_5;
wire [7:0] nScanOut1733;
wire [7:0] nOut27_6;
wire [7:0] nScanOut1734;
wire [7:0] nOut27_7;
wire [7:0] nScanOut1735;
wire [7:0] nOut27_8;
wire [7:0] nScanOut1736;
wire [7:0] nOut27_9;
wire [7:0] nScanOut1737;
wire [7:0] nOut27_10;
wire [7:0] nScanOut1738;
wire [7:0] nOut27_11;
wire [7:0] nScanOut1739;
wire [7:0] nOut27_12;
wire [7:0] nScanOut1740;
wire [7:0] nOut27_13;
wire [7:0] nScanOut1741;
wire [7:0] nOut27_14;
wire [7:0] nScanOut1742;
wire [7:0] nOut27_15;
wire [7:0] nScanOut1743;
wire [7:0] nOut27_16;
wire [7:0] nScanOut1744;
wire [7:0] nOut27_17;
wire [7:0] nScanOut1745;
wire [7:0] nOut27_18;
wire [7:0] nScanOut1746;
wire [7:0] nOut27_19;
wire [7:0] nScanOut1747;
wire [7:0] nOut27_20;
wire [7:0] nScanOut1748;
wire [7:0] nOut27_21;
wire [7:0] nScanOut1749;
wire [7:0] nOut27_22;
wire [7:0] nScanOut1750;
wire [7:0] nOut27_23;
wire [7:0] nScanOut1751;
wire [7:0] nOut27_24;
wire [7:0] nScanOut1752;
wire [7:0] nOut27_25;
wire [7:0] nScanOut1753;
wire [7:0] nOut27_26;
wire [7:0] nScanOut1754;
wire [7:0] nOut27_27;
wire [7:0] nScanOut1755;
wire [7:0] nOut27_28;
wire [7:0] nScanOut1756;
wire [7:0] nOut27_29;
wire [7:0] nScanOut1757;
wire [7:0] nOut27_30;
wire [7:0] nScanOut1758;
wire [7:0] nOut27_31;
wire [7:0] nScanOut1759;
wire [7:0] nOut27_32;
wire [7:0] nScanOut1760;
wire [7:0] nOut27_33;
wire [7:0] nScanOut1761;
wire [7:0] nOut27_34;
wire [7:0] nScanOut1762;
wire [7:0] nOut27_35;
wire [7:0] nScanOut1763;
wire [7:0] nOut27_36;
wire [7:0] nScanOut1764;
wire [7:0] nOut27_37;
wire [7:0] nScanOut1765;
wire [7:0] nOut27_38;
wire [7:0] nScanOut1766;
wire [7:0] nOut27_39;
wire [7:0] nScanOut1767;
wire [7:0] nOut27_40;
wire [7:0] nScanOut1768;
wire [7:0] nOut27_41;
wire [7:0] nScanOut1769;
wire [7:0] nOut27_42;
wire [7:0] nScanOut1770;
wire [7:0] nOut27_43;
wire [7:0] nScanOut1771;
wire [7:0] nOut27_44;
wire [7:0] nScanOut1772;
wire [7:0] nOut27_45;
wire [7:0] nScanOut1773;
wire [7:0] nOut27_46;
wire [7:0] nScanOut1774;
wire [7:0] nOut27_47;
wire [7:0] nScanOut1775;
wire [7:0] nOut27_48;
wire [7:0] nScanOut1776;
wire [7:0] nOut27_49;
wire [7:0] nScanOut1777;
wire [7:0] nOut27_50;
wire [7:0] nScanOut1778;
wire [7:0] nOut27_51;
wire [7:0] nScanOut1779;
wire [7:0] nOut27_52;
wire [7:0] nScanOut1780;
wire [7:0] nOut27_53;
wire [7:0] nScanOut1781;
wire [7:0] nOut27_54;
wire [7:0] nScanOut1782;
wire [7:0] nOut27_55;
wire [7:0] nScanOut1783;
wire [7:0] nOut27_56;
wire [7:0] nScanOut1784;
wire [7:0] nOut27_57;
wire [7:0] nScanOut1785;
wire [7:0] nOut27_58;
wire [7:0] nScanOut1786;
wire [7:0] nOut27_59;
wire [7:0] nScanOut1787;
wire [7:0] nOut27_60;
wire [7:0] nScanOut1788;
wire [7:0] nOut27_61;
wire [7:0] nScanOut1789;
wire [7:0] nOut27_62;
wire [7:0] nScanOut1790;
wire [7:0] nOut27_63;
wire [7:0] nScanOut1791;
wire [7:0] nOut28_0;
wire [7:0] nScanOut1792;
wire [7:0] nOut28_1;
wire [7:0] nScanOut1793;
wire [7:0] nOut28_2;
wire [7:0] nScanOut1794;
wire [7:0] nOut28_3;
wire [7:0] nScanOut1795;
wire [7:0] nOut28_4;
wire [7:0] nScanOut1796;
wire [7:0] nOut28_5;
wire [7:0] nScanOut1797;
wire [7:0] nOut28_6;
wire [7:0] nScanOut1798;
wire [7:0] nOut28_7;
wire [7:0] nScanOut1799;
wire [7:0] nOut28_8;
wire [7:0] nScanOut1800;
wire [7:0] nOut28_9;
wire [7:0] nScanOut1801;
wire [7:0] nOut28_10;
wire [7:0] nScanOut1802;
wire [7:0] nOut28_11;
wire [7:0] nScanOut1803;
wire [7:0] nOut28_12;
wire [7:0] nScanOut1804;
wire [7:0] nOut28_13;
wire [7:0] nScanOut1805;
wire [7:0] nOut28_14;
wire [7:0] nScanOut1806;
wire [7:0] nOut28_15;
wire [7:0] nScanOut1807;
wire [7:0] nOut28_16;
wire [7:0] nScanOut1808;
wire [7:0] nOut28_17;
wire [7:0] nScanOut1809;
wire [7:0] nOut28_18;
wire [7:0] nScanOut1810;
wire [7:0] nOut28_19;
wire [7:0] nScanOut1811;
wire [7:0] nOut28_20;
wire [7:0] nScanOut1812;
wire [7:0] nOut28_21;
wire [7:0] nScanOut1813;
wire [7:0] nOut28_22;
wire [7:0] nScanOut1814;
wire [7:0] nOut28_23;
wire [7:0] nScanOut1815;
wire [7:0] nOut28_24;
wire [7:0] nScanOut1816;
wire [7:0] nOut28_25;
wire [7:0] nScanOut1817;
wire [7:0] nOut28_26;
wire [7:0] nScanOut1818;
wire [7:0] nOut28_27;
wire [7:0] nScanOut1819;
wire [7:0] nOut28_28;
wire [7:0] nScanOut1820;
wire [7:0] nOut28_29;
wire [7:0] nScanOut1821;
wire [7:0] nOut28_30;
wire [7:0] nScanOut1822;
wire [7:0] nOut28_31;
wire [7:0] nScanOut1823;
wire [7:0] nOut28_32;
wire [7:0] nScanOut1824;
wire [7:0] nOut28_33;
wire [7:0] nScanOut1825;
wire [7:0] nOut28_34;
wire [7:0] nScanOut1826;
wire [7:0] nOut28_35;
wire [7:0] nScanOut1827;
wire [7:0] nOut28_36;
wire [7:0] nScanOut1828;
wire [7:0] nOut28_37;
wire [7:0] nScanOut1829;
wire [7:0] nOut28_38;
wire [7:0] nScanOut1830;
wire [7:0] nOut28_39;
wire [7:0] nScanOut1831;
wire [7:0] nOut28_40;
wire [7:0] nScanOut1832;
wire [7:0] nOut28_41;
wire [7:0] nScanOut1833;
wire [7:0] nOut28_42;
wire [7:0] nScanOut1834;
wire [7:0] nOut28_43;
wire [7:0] nScanOut1835;
wire [7:0] nOut28_44;
wire [7:0] nScanOut1836;
wire [7:0] nOut28_45;
wire [7:0] nScanOut1837;
wire [7:0] nOut28_46;
wire [7:0] nScanOut1838;
wire [7:0] nOut28_47;
wire [7:0] nScanOut1839;
wire [7:0] nOut28_48;
wire [7:0] nScanOut1840;
wire [7:0] nOut28_49;
wire [7:0] nScanOut1841;
wire [7:0] nOut28_50;
wire [7:0] nScanOut1842;
wire [7:0] nOut28_51;
wire [7:0] nScanOut1843;
wire [7:0] nOut28_52;
wire [7:0] nScanOut1844;
wire [7:0] nOut28_53;
wire [7:0] nScanOut1845;
wire [7:0] nOut28_54;
wire [7:0] nScanOut1846;
wire [7:0] nOut28_55;
wire [7:0] nScanOut1847;
wire [7:0] nOut28_56;
wire [7:0] nScanOut1848;
wire [7:0] nOut28_57;
wire [7:0] nScanOut1849;
wire [7:0] nOut28_58;
wire [7:0] nScanOut1850;
wire [7:0] nOut28_59;
wire [7:0] nScanOut1851;
wire [7:0] nOut28_60;
wire [7:0] nScanOut1852;
wire [7:0] nOut28_61;
wire [7:0] nScanOut1853;
wire [7:0] nOut28_62;
wire [7:0] nScanOut1854;
wire [7:0] nOut28_63;
wire [7:0] nScanOut1855;
wire [7:0] nOut29_0;
wire [7:0] nScanOut1856;
wire [7:0] nOut29_1;
wire [7:0] nScanOut1857;
wire [7:0] nOut29_2;
wire [7:0] nScanOut1858;
wire [7:0] nOut29_3;
wire [7:0] nScanOut1859;
wire [7:0] nOut29_4;
wire [7:0] nScanOut1860;
wire [7:0] nOut29_5;
wire [7:0] nScanOut1861;
wire [7:0] nOut29_6;
wire [7:0] nScanOut1862;
wire [7:0] nOut29_7;
wire [7:0] nScanOut1863;
wire [7:0] nOut29_8;
wire [7:0] nScanOut1864;
wire [7:0] nOut29_9;
wire [7:0] nScanOut1865;
wire [7:0] nOut29_10;
wire [7:0] nScanOut1866;
wire [7:0] nOut29_11;
wire [7:0] nScanOut1867;
wire [7:0] nOut29_12;
wire [7:0] nScanOut1868;
wire [7:0] nOut29_13;
wire [7:0] nScanOut1869;
wire [7:0] nOut29_14;
wire [7:0] nScanOut1870;
wire [7:0] nOut29_15;
wire [7:0] nScanOut1871;
wire [7:0] nOut29_16;
wire [7:0] nScanOut1872;
wire [7:0] nOut29_17;
wire [7:0] nScanOut1873;
wire [7:0] nOut29_18;
wire [7:0] nScanOut1874;
wire [7:0] nOut29_19;
wire [7:0] nScanOut1875;
wire [7:0] nOut29_20;
wire [7:0] nScanOut1876;
wire [7:0] nOut29_21;
wire [7:0] nScanOut1877;
wire [7:0] nOut29_22;
wire [7:0] nScanOut1878;
wire [7:0] nOut29_23;
wire [7:0] nScanOut1879;
wire [7:0] nOut29_24;
wire [7:0] nScanOut1880;
wire [7:0] nOut29_25;
wire [7:0] nScanOut1881;
wire [7:0] nOut29_26;
wire [7:0] nScanOut1882;
wire [7:0] nOut29_27;
wire [7:0] nScanOut1883;
wire [7:0] nOut29_28;
wire [7:0] nScanOut1884;
wire [7:0] nOut29_29;
wire [7:0] nScanOut1885;
wire [7:0] nOut29_30;
wire [7:0] nScanOut1886;
wire [7:0] nOut29_31;
wire [7:0] nScanOut1887;
wire [7:0] nOut29_32;
wire [7:0] nScanOut1888;
wire [7:0] nOut29_33;
wire [7:0] nScanOut1889;
wire [7:0] nOut29_34;
wire [7:0] nScanOut1890;
wire [7:0] nOut29_35;
wire [7:0] nScanOut1891;
wire [7:0] nOut29_36;
wire [7:0] nScanOut1892;
wire [7:0] nOut29_37;
wire [7:0] nScanOut1893;
wire [7:0] nOut29_38;
wire [7:0] nScanOut1894;
wire [7:0] nOut29_39;
wire [7:0] nScanOut1895;
wire [7:0] nOut29_40;
wire [7:0] nScanOut1896;
wire [7:0] nOut29_41;
wire [7:0] nScanOut1897;
wire [7:0] nOut29_42;
wire [7:0] nScanOut1898;
wire [7:0] nOut29_43;
wire [7:0] nScanOut1899;
wire [7:0] nOut29_44;
wire [7:0] nScanOut1900;
wire [7:0] nOut29_45;
wire [7:0] nScanOut1901;
wire [7:0] nOut29_46;
wire [7:0] nScanOut1902;
wire [7:0] nOut29_47;
wire [7:0] nScanOut1903;
wire [7:0] nOut29_48;
wire [7:0] nScanOut1904;
wire [7:0] nOut29_49;
wire [7:0] nScanOut1905;
wire [7:0] nOut29_50;
wire [7:0] nScanOut1906;
wire [7:0] nOut29_51;
wire [7:0] nScanOut1907;
wire [7:0] nOut29_52;
wire [7:0] nScanOut1908;
wire [7:0] nOut29_53;
wire [7:0] nScanOut1909;
wire [7:0] nOut29_54;
wire [7:0] nScanOut1910;
wire [7:0] nOut29_55;
wire [7:0] nScanOut1911;
wire [7:0] nOut29_56;
wire [7:0] nScanOut1912;
wire [7:0] nOut29_57;
wire [7:0] nScanOut1913;
wire [7:0] nOut29_58;
wire [7:0] nScanOut1914;
wire [7:0] nOut29_59;
wire [7:0] nScanOut1915;
wire [7:0] nOut29_60;
wire [7:0] nScanOut1916;
wire [7:0] nOut29_61;
wire [7:0] nScanOut1917;
wire [7:0] nOut29_62;
wire [7:0] nScanOut1918;
wire [7:0] nOut29_63;
wire [7:0] nScanOut1919;
wire [7:0] nOut30_0;
wire [7:0] nScanOut1920;
wire [7:0] nOut30_1;
wire [7:0] nScanOut1921;
wire [7:0] nOut30_2;
wire [7:0] nScanOut1922;
wire [7:0] nOut30_3;
wire [7:0] nScanOut1923;
wire [7:0] nOut30_4;
wire [7:0] nScanOut1924;
wire [7:0] nOut30_5;
wire [7:0] nScanOut1925;
wire [7:0] nOut30_6;
wire [7:0] nScanOut1926;
wire [7:0] nOut30_7;
wire [7:0] nScanOut1927;
wire [7:0] nOut30_8;
wire [7:0] nScanOut1928;
wire [7:0] nOut30_9;
wire [7:0] nScanOut1929;
wire [7:0] nOut30_10;
wire [7:0] nScanOut1930;
wire [7:0] nOut30_11;
wire [7:0] nScanOut1931;
wire [7:0] nOut30_12;
wire [7:0] nScanOut1932;
wire [7:0] nOut30_13;
wire [7:0] nScanOut1933;
wire [7:0] nOut30_14;
wire [7:0] nScanOut1934;
wire [7:0] nOut30_15;
wire [7:0] nScanOut1935;
wire [7:0] nOut30_16;
wire [7:0] nScanOut1936;
wire [7:0] nOut30_17;
wire [7:0] nScanOut1937;
wire [7:0] nOut30_18;
wire [7:0] nScanOut1938;
wire [7:0] nOut30_19;
wire [7:0] nScanOut1939;
wire [7:0] nOut30_20;
wire [7:0] nScanOut1940;
wire [7:0] nOut30_21;
wire [7:0] nScanOut1941;
wire [7:0] nOut30_22;
wire [7:0] nScanOut1942;
wire [7:0] nOut30_23;
wire [7:0] nScanOut1943;
wire [7:0] nOut30_24;
wire [7:0] nScanOut1944;
wire [7:0] nOut30_25;
wire [7:0] nScanOut1945;
wire [7:0] nOut30_26;
wire [7:0] nScanOut1946;
wire [7:0] nOut30_27;
wire [7:0] nScanOut1947;
wire [7:0] nOut30_28;
wire [7:0] nScanOut1948;
wire [7:0] nOut30_29;
wire [7:0] nScanOut1949;
wire [7:0] nOut30_30;
wire [7:0] nScanOut1950;
wire [7:0] nOut30_31;
wire [7:0] nScanOut1951;
wire [7:0] nOut30_32;
wire [7:0] nScanOut1952;
wire [7:0] nOut30_33;
wire [7:0] nScanOut1953;
wire [7:0] nOut30_34;
wire [7:0] nScanOut1954;
wire [7:0] nOut30_35;
wire [7:0] nScanOut1955;
wire [7:0] nOut30_36;
wire [7:0] nScanOut1956;
wire [7:0] nOut30_37;
wire [7:0] nScanOut1957;
wire [7:0] nOut30_38;
wire [7:0] nScanOut1958;
wire [7:0] nOut30_39;
wire [7:0] nScanOut1959;
wire [7:0] nOut30_40;
wire [7:0] nScanOut1960;
wire [7:0] nOut30_41;
wire [7:0] nScanOut1961;
wire [7:0] nOut30_42;
wire [7:0] nScanOut1962;
wire [7:0] nOut30_43;
wire [7:0] nScanOut1963;
wire [7:0] nOut30_44;
wire [7:0] nScanOut1964;
wire [7:0] nOut30_45;
wire [7:0] nScanOut1965;
wire [7:0] nOut30_46;
wire [7:0] nScanOut1966;
wire [7:0] nOut30_47;
wire [7:0] nScanOut1967;
wire [7:0] nOut30_48;
wire [7:0] nScanOut1968;
wire [7:0] nOut30_49;
wire [7:0] nScanOut1969;
wire [7:0] nOut30_50;
wire [7:0] nScanOut1970;
wire [7:0] nOut30_51;
wire [7:0] nScanOut1971;
wire [7:0] nOut30_52;
wire [7:0] nScanOut1972;
wire [7:0] nOut30_53;
wire [7:0] nScanOut1973;
wire [7:0] nOut30_54;
wire [7:0] nScanOut1974;
wire [7:0] nOut30_55;
wire [7:0] nScanOut1975;
wire [7:0] nOut30_56;
wire [7:0] nScanOut1976;
wire [7:0] nOut30_57;
wire [7:0] nScanOut1977;
wire [7:0] nOut30_58;
wire [7:0] nScanOut1978;
wire [7:0] nOut30_59;
wire [7:0] nScanOut1979;
wire [7:0] nOut30_60;
wire [7:0] nScanOut1980;
wire [7:0] nOut30_61;
wire [7:0] nScanOut1981;
wire [7:0] nOut30_62;
wire [7:0] nScanOut1982;
wire [7:0] nOut30_63;
wire [7:0] nScanOut1983;
wire [7:0] nOut31_0;
wire [7:0] nScanOut1984;
wire [7:0] nOut31_1;
wire [7:0] nScanOut1985;
wire [7:0] nOut31_2;
wire [7:0] nScanOut1986;
wire [7:0] nOut31_3;
wire [7:0] nScanOut1987;
wire [7:0] nOut31_4;
wire [7:0] nScanOut1988;
wire [7:0] nOut31_5;
wire [7:0] nScanOut1989;
wire [7:0] nOut31_6;
wire [7:0] nScanOut1990;
wire [7:0] nOut31_7;
wire [7:0] nScanOut1991;
wire [7:0] nOut31_8;
wire [7:0] nScanOut1992;
wire [7:0] nOut31_9;
wire [7:0] nScanOut1993;
wire [7:0] nOut31_10;
wire [7:0] nScanOut1994;
wire [7:0] nOut31_11;
wire [7:0] nScanOut1995;
wire [7:0] nOut31_12;
wire [7:0] nScanOut1996;
wire [7:0] nOut31_13;
wire [7:0] nScanOut1997;
wire [7:0] nOut31_14;
wire [7:0] nScanOut1998;
wire [7:0] nOut31_15;
wire [7:0] nScanOut1999;
wire [7:0] nOut31_16;
wire [7:0] nScanOut2000;
wire [7:0] nOut31_17;
wire [7:0] nScanOut2001;
wire [7:0] nOut31_18;
wire [7:0] nScanOut2002;
wire [7:0] nOut31_19;
wire [7:0] nScanOut2003;
wire [7:0] nOut31_20;
wire [7:0] nScanOut2004;
wire [7:0] nOut31_21;
wire [7:0] nScanOut2005;
wire [7:0] nOut31_22;
wire [7:0] nScanOut2006;
wire [7:0] nOut31_23;
wire [7:0] nScanOut2007;
wire [7:0] nOut31_24;
wire [7:0] nScanOut2008;
wire [7:0] nOut31_25;
wire [7:0] nScanOut2009;
wire [7:0] nOut31_26;
wire [7:0] nScanOut2010;
wire [7:0] nOut31_27;
wire [7:0] nScanOut2011;
wire [7:0] nOut31_28;
wire [7:0] nScanOut2012;
wire [7:0] nOut31_29;
wire [7:0] nScanOut2013;
wire [7:0] nOut31_30;
wire [7:0] nScanOut2014;
wire [7:0] nOut31_31;
wire [7:0] nScanOut2015;
wire [7:0] nOut31_32;
wire [7:0] nScanOut2016;
wire [7:0] nOut31_33;
wire [7:0] nScanOut2017;
wire [7:0] nOut31_34;
wire [7:0] nScanOut2018;
wire [7:0] nOut31_35;
wire [7:0] nScanOut2019;
wire [7:0] nOut31_36;
wire [7:0] nScanOut2020;
wire [7:0] nOut31_37;
wire [7:0] nScanOut2021;
wire [7:0] nOut31_38;
wire [7:0] nScanOut2022;
wire [7:0] nOut31_39;
wire [7:0] nScanOut2023;
wire [7:0] nOut31_40;
wire [7:0] nScanOut2024;
wire [7:0] nOut31_41;
wire [7:0] nScanOut2025;
wire [7:0] nOut31_42;
wire [7:0] nScanOut2026;
wire [7:0] nOut31_43;
wire [7:0] nScanOut2027;
wire [7:0] nOut31_44;
wire [7:0] nScanOut2028;
wire [7:0] nOut31_45;
wire [7:0] nScanOut2029;
wire [7:0] nOut31_46;
wire [7:0] nScanOut2030;
wire [7:0] nOut31_47;
wire [7:0] nScanOut2031;
wire [7:0] nOut31_48;
wire [7:0] nScanOut2032;
wire [7:0] nOut31_49;
wire [7:0] nScanOut2033;
wire [7:0] nOut31_50;
wire [7:0] nScanOut2034;
wire [7:0] nOut31_51;
wire [7:0] nScanOut2035;
wire [7:0] nOut31_52;
wire [7:0] nScanOut2036;
wire [7:0] nOut31_53;
wire [7:0] nScanOut2037;
wire [7:0] nOut31_54;
wire [7:0] nScanOut2038;
wire [7:0] nOut31_55;
wire [7:0] nScanOut2039;
wire [7:0] nOut31_56;
wire [7:0] nScanOut2040;
wire [7:0] nOut31_57;
wire [7:0] nScanOut2041;
wire [7:0] nOut31_58;
wire [7:0] nScanOut2042;
wire [7:0] nOut31_59;
wire [7:0] nScanOut2043;
wire [7:0] nOut31_60;
wire [7:0] nScanOut2044;
wire [7:0] nOut31_61;
wire [7:0] nScanOut2045;
wire [7:0] nOut31_62;
wire [7:0] nScanOut2046;
wire [7:0] nOut31_63;
wire [7:0] nScanOut2047;
wire [0:0] nEnable;
wire [0:0] nScanEnable;
wire [7:0] nScanOut2048;
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_0), .ScanIn(nScanOut1), .ScanOut(nScanOut0), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_1), .ScanIn(nScanOut2), .ScanOut(nScanOut1), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_2), .ScanIn(nScanOut3), .ScanOut(nScanOut2), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_3), .ScanIn(nScanOut4), .ScanOut(nScanOut3), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_4), .ScanIn(nScanOut5), .ScanOut(nScanOut4), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_5), .ScanIn(nScanOut6), .ScanOut(nScanOut5), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_6), .ScanIn(nScanOut7), .ScanOut(nScanOut6), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_7), .ScanIn(nScanOut8), .ScanOut(nScanOut7), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_8), .ScanIn(nScanOut9), .ScanOut(nScanOut8), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_9), .ScanIn(nScanOut10), .ScanOut(nScanOut9), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_10), .ScanIn(nScanOut11), .ScanOut(nScanOut10), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_11), .ScanIn(nScanOut12), .ScanOut(nScanOut11), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_12), .ScanIn(nScanOut13), .ScanOut(nScanOut12), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_13), .ScanIn(nScanOut14), .ScanOut(nScanOut13), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_14), .ScanIn(nScanOut15), .ScanOut(nScanOut14), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_15), .ScanIn(nScanOut16), .ScanOut(nScanOut15), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_16), .ScanIn(nScanOut17), .ScanOut(nScanOut16), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_17), .ScanIn(nScanOut18), .ScanOut(nScanOut17), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_18), .ScanIn(nScanOut19), .ScanOut(nScanOut18), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_19), .ScanIn(nScanOut20), .ScanOut(nScanOut19), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_20), .ScanIn(nScanOut21), .ScanOut(nScanOut20), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_21), .ScanIn(nScanOut22), .ScanOut(nScanOut21), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_22), .ScanIn(nScanOut23), .ScanOut(nScanOut22), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_23), .ScanIn(nScanOut24), .ScanOut(nScanOut23), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_24), .ScanIn(nScanOut25), .ScanOut(nScanOut24), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_25), .ScanIn(nScanOut26), .ScanOut(nScanOut25), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_26), .ScanIn(nScanOut27), .ScanOut(nScanOut26), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_27), .ScanIn(nScanOut28), .ScanOut(nScanOut27), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_28), .ScanIn(nScanOut29), .ScanOut(nScanOut28), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_29), .ScanIn(nScanOut30), .ScanOut(nScanOut29), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_30), .ScanIn(nScanOut31), .ScanOut(nScanOut30), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_31), .ScanIn(nScanOut32), .ScanOut(nScanOut31), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_32), .ScanIn(nScanOut33), .ScanOut(nScanOut32), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_33), .ScanIn(nScanOut34), .ScanOut(nScanOut33), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_34), .ScanIn(nScanOut35), .ScanOut(nScanOut34), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_35), .ScanIn(nScanOut36), .ScanOut(nScanOut35), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_36), .ScanIn(nScanOut37), .ScanOut(nScanOut36), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_37), .ScanIn(nScanOut38), .ScanOut(nScanOut37), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_38), .ScanIn(nScanOut39), .ScanOut(nScanOut38), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_39), .ScanIn(nScanOut40), .ScanOut(nScanOut39), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_40), .ScanIn(nScanOut41), .ScanOut(nScanOut40), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_41), .ScanIn(nScanOut42), .ScanOut(nScanOut41), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_42), .ScanIn(nScanOut43), .ScanOut(nScanOut42), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_43), .ScanIn(nScanOut44), .ScanOut(nScanOut43), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_44), .ScanIn(nScanOut45), .ScanOut(nScanOut44), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_45), .ScanIn(nScanOut46), .ScanOut(nScanOut45), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_46), .ScanIn(nScanOut47), .ScanOut(nScanOut46), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_47), .ScanIn(nScanOut48), .ScanOut(nScanOut47), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_48), .ScanIn(nScanOut49), .ScanOut(nScanOut48), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_49), .ScanIn(nScanOut50), .ScanOut(nScanOut49), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_50), .ScanIn(nScanOut51), .ScanOut(nScanOut50), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_51), .ScanIn(nScanOut52), .ScanOut(nScanOut51), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_52), .ScanIn(nScanOut53), .ScanOut(nScanOut52), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_53), .ScanIn(nScanOut54), .ScanOut(nScanOut53), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_54), .ScanIn(nScanOut55), .ScanOut(nScanOut54), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_55), .ScanIn(nScanOut56), .ScanOut(nScanOut55), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_56), .ScanIn(nScanOut57), .ScanOut(nScanOut56), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_57), .ScanIn(nScanOut58), .ScanOut(nScanOut57), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_58), .ScanIn(nScanOut59), .ScanOut(nScanOut58), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_59), .ScanIn(nScanOut60), .ScanOut(nScanOut59), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_60), .ScanIn(nScanOut61), .ScanOut(nScanOut60), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_61), .ScanIn(nScanOut62), .ScanOut(nScanOut61), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_62), .ScanIn(nScanOut63), .ScanOut(nScanOut62), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_63), .ScanIn(nScanOut64), .ScanOut(nScanOut63), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_0), .ScanIn(nScanOut65), .ScanOut(nScanOut64), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_1), .NorthIn(nOut1_0), .SouthIn(nOut1_2), .EastIn(nOut2_1), .WestIn(nOut0_1), .ScanIn(nScanOut66), .ScanOut(nScanOut65), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_2), .NorthIn(nOut1_1), .SouthIn(nOut1_3), .EastIn(nOut2_2), .WestIn(nOut0_2), .ScanIn(nScanOut67), .ScanOut(nScanOut66), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_3), .NorthIn(nOut1_2), .SouthIn(nOut1_4), .EastIn(nOut2_3), .WestIn(nOut0_3), .ScanIn(nScanOut68), .ScanOut(nScanOut67), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_4), .NorthIn(nOut1_3), .SouthIn(nOut1_5), .EastIn(nOut2_4), .WestIn(nOut0_4), .ScanIn(nScanOut69), .ScanOut(nScanOut68), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_5), .NorthIn(nOut1_4), .SouthIn(nOut1_6), .EastIn(nOut2_5), .WestIn(nOut0_5), .ScanIn(nScanOut70), .ScanOut(nScanOut69), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_6), .NorthIn(nOut1_5), .SouthIn(nOut1_7), .EastIn(nOut2_6), .WestIn(nOut0_6), .ScanIn(nScanOut71), .ScanOut(nScanOut70), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_7), .NorthIn(nOut1_6), .SouthIn(nOut1_8), .EastIn(nOut2_7), .WestIn(nOut0_7), .ScanIn(nScanOut72), .ScanOut(nScanOut71), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_8), .NorthIn(nOut1_7), .SouthIn(nOut1_9), .EastIn(nOut2_8), .WestIn(nOut0_8), .ScanIn(nScanOut73), .ScanOut(nScanOut72), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_9), .NorthIn(nOut1_8), .SouthIn(nOut1_10), .EastIn(nOut2_9), .WestIn(nOut0_9), .ScanIn(nScanOut74), .ScanOut(nScanOut73), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_10), .NorthIn(nOut1_9), .SouthIn(nOut1_11), .EastIn(nOut2_10), .WestIn(nOut0_10), .ScanIn(nScanOut75), .ScanOut(nScanOut74), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_11), .NorthIn(nOut1_10), .SouthIn(nOut1_12), .EastIn(nOut2_11), .WestIn(nOut0_11), .ScanIn(nScanOut76), .ScanOut(nScanOut75), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_12), .NorthIn(nOut1_11), .SouthIn(nOut1_13), .EastIn(nOut2_12), .WestIn(nOut0_12), .ScanIn(nScanOut77), .ScanOut(nScanOut76), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_13), .NorthIn(nOut1_12), .SouthIn(nOut1_14), .EastIn(nOut2_13), .WestIn(nOut0_13), .ScanIn(nScanOut78), .ScanOut(nScanOut77), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_14), .NorthIn(nOut1_13), .SouthIn(nOut1_15), .EastIn(nOut2_14), .WestIn(nOut0_14), .ScanIn(nScanOut79), .ScanOut(nScanOut78), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_15), .NorthIn(nOut1_14), .SouthIn(nOut1_16), .EastIn(nOut2_15), .WestIn(nOut0_15), .ScanIn(nScanOut80), .ScanOut(nScanOut79), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_16), .NorthIn(nOut1_15), .SouthIn(nOut1_17), .EastIn(nOut2_16), .WestIn(nOut0_16), .ScanIn(nScanOut81), .ScanOut(nScanOut80), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_17), .NorthIn(nOut1_16), .SouthIn(nOut1_18), .EastIn(nOut2_17), .WestIn(nOut0_17), .ScanIn(nScanOut82), .ScanOut(nScanOut81), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_18), .NorthIn(nOut1_17), .SouthIn(nOut1_19), .EastIn(nOut2_18), .WestIn(nOut0_18), .ScanIn(nScanOut83), .ScanOut(nScanOut82), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_19), .NorthIn(nOut1_18), .SouthIn(nOut1_20), .EastIn(nOut2_19), .WestIn(nOut0_19), .ScanIn(nScanOut84), .ScanOut(nScanOut83), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_20), .NorthIn(nOut1_19), .SouthIn(nOut1_21), .EastIn(nOut2_20), .WestIn(nOut0_20), .ScanIn(nScanOut85), .ScanOut(nScanOut84), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_21), .NorthIn(nOut1_20), .SouthIn(nOut1_22), .EastIn(nOut2_21), .WestIn(nOut0_21), .ScanIn(nScanOut86), .ScanOut(nScanOut85), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_22), .NorthIn(nOut1_21), .SouthIn(nOut1_23), .EastIn(nOut2_22), .WestIn(nOut0_22), .ScanIn(nScanOut87), .ScanOut(nScanOut86), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_23), .NorthIn(nOut1_22), .SouthIn(nOut1_24), .EastIn(nOut2_23), .WestIn(nOut0_23), .ScanIn(nScanOut88), .ScanOut(nScanOut87), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_24), .NorthIn(nOut1_23), .SouthIn(nOut1_25), .EastIn(nOut2_24), .WestIn(nOut0_24), .ScanIn(nScanOut89), .ScanOut(nScanOut88), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_25), .NorthIn(nOut1_24), .SouthIn(nOut1_26), .EastIn(nOut2_25), .WestIn(nOut0_25), .ScanIn(nScanOut90), .ScanOut(nScanOut89), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_26), .NorthIn(nOut1_25), .SouthIn(nOut1_27), .EastIn(nOut2_26), .WestIn(nOut0_26), .ScanIn(nScanOut91), .ScanOut(nScanOut90), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_27), .NorthIn(nOut1_26), .SouthIn(nOut1_28), .EastIn(nOut2_27), .WestIn(nOut0_27), .ScanIn(nScanOut92), .ScanOut(nScanOut91), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_28), .NorthIn(nOut1_27), .SouthIn(nOut1_29), .EastIn(nOut2_28), .WestIn(nOut0_28), .ScanIn(nScanOut93), .ScanOut(nScanOut92), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_29), .NorthIn(nOut1_28), .SouthIn(nOut1_30), .EastIn(nOut2_29), .WestIn(nOut0_29), .ScanIn(nScanOut94), .ScanOut(nScanOut93), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_30), .NorthIn(nOut1_29), .SouthIn(nOut1_31), .EastIn(nOut2_30), .WestIn(nOut0_30), .ScanIn(nScanOut95), .ScanOut(nScanOut94), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_31), .NorthIn(nOut1_30), .SouthIn(nOut1_32), .EastIn(nOut2_31), .WestIn(nOut0_31), .ScanIn(nScanOut96), .ScanOut(nScanOut95), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_32), .NorthIn(nOut1_31), .SouthIn(nOut1_33), .EastIn(nOut2_32), .WestIn(nOut0_32), .ScanIn(nScanOut97), .ScanOut(nScanOut96), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_33), .NorthIn(nOut1_32), .SouthIn(nOut1_34), .EastIn(nOut2_33), .WestIn(nOut0_33), .ScanIn(nScanOut98), .ScanOut(nScanOut97), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_34), .NorthIn(nOut1_33), .SouthIn(nOut1_35), .EastIn(nOut2_34), .WestIn(nOut0_34), .ScanIn(nScanOut99), .ScanOut(nScanOut98), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_35), .NorthIn(nOut1_34), .SouthIn(nOut1_36), .EastIn(nOut2_35), .WestIn(nOut0_35), .ScanIn(nScanOut100), .ScanOut(nScanOut99), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_36), .NorthIn(nOut1_35), .SouthIn(nOut1_37), .EastIn(nOut2_36), .WestIn(nOut0_36), .ScanIn(nScanOut101), .ScanOut(nScanOut100), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_37), .NorthIn(nOut1_36), .SouthIn(nOut1_38), .EastIn(nOut2_37), .WestIn(nOut0_37), .ScanIn(nScanOut102), .ScanOut(nScanOut101), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_38), .NorthIn(nOut1_37), .SouthIn(nOut1_39), .EastIn(nOut2_38), .WestIn(nOut0_38), .ScanIn(nScanOut103), .ScanOut(nScanOut102), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_39), .NorthIn(nOut1_38), .SouthIn(nOut1_40), .EastIn(nOut2_39), .WestIn(nOut0_39), .ScanIn(nScanOut104), .ScanOut(nScanOut103), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_40), .NorthIn(nOut1_39), .SouthIn(nOut1_41), .EastIn(nOut2_40), .WestIn(nOut0_40), .ScanIn(nScanOut105), .ScanOut(nScanOut104), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_41), .NorthIn(nOut1_40), .SouthIn(nOut1_42), .EastIn(nOut2_41), .WestIn(nOut0_41), .ScanIn(nScanOut106), .ScanOut(nScanOut105), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_42), .NorthIn(nOut1_41), .SouthIn(nOut1_43), .EastIn(nOut2_42), .WestIn(nOut0_42), .ScanIn(nScanOut107), .ScanOut(nScanOut106), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_43), .NorthIn(nOut1_42), .SouthIn(nOut1_44), .EastIn(nOut2_43), .WestIn(nOut0_43), .ScanIn(nScanOut108), .ScanOut(nScanOut107), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_44), .NorthIn(nOut1_43), .SouthIn(nOut1_45), .EastIn(nOut2_44), .WestIn(nOut0_44), .ScanIn(nScanOut109), .ScanOut(nScanOut108), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_45), .NorthIn(nOut1_44), .SouthIn(nOut1_46), .EastIn(nOut2_45), .WestIn(nOut0_45), .ScanIn(nScanOut110), .ScanOut(nScanOut109), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_46), .NorthIn(nOut1_45), .SouthIn(nOut1_47), .EastIn(nOut2_46), .WestIn(nOut0_46), .ScanIn(nScanOut111), .ScanOut(nScanOut110), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_47), .NorthIn(nOut1_46), .SouthIn(nOut1_48), .EastIn(nOut2_47), .WestIn(nOut0_47), .ScanIn(nScanOut112), .ScanOut(nScanOut111), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_48), .NorthIn(nOut1_47), .SouthIn(nOut1_49), .EastIn(nOut2_48), .WestIn(nOut0_48), .ScanIn(nScanOut113), .ScanOut(nScanOut112), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_49), .NorthIn(nOut1_48), .SouthIn(nOut1_50), .EastIn(nOut2_49), .WestIn(nOut0_49), .ScanIn(nScanOut114), .ScanOut(nScanOut113), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_50), .NorthIn(nOut1_49), .SouthIn(nOut1_51), .EastIn(nOut2_50), .WestIn(nOut0_50), .ScanIn(nScanOut115), .ScanOut(nScanOut114), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_51), .NorthIn(nOut1_50), .SouthIn(nOut1_52), .EastIn(nOut2_51), .WestIn(nOut0_51), .ScanIn(nScanOut116), .ScanOut(nScanOut115), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_52), .NorthIn(nOut1_51), .SouthIn(nOut1_53), .EastIn(nOut2_52), .WestIn(nOut0_52), .ScanIn(nScanOut117), .ScanOut(nScanOut116), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_53), .NorthIn(nOut1_52), .SouthIn(nOut1_54), .EastIn(nOut2_53), .WestIn(nOut0_53), .ScanIn(nScanOut118), .ScanOut(nScanOut117), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_54), .NorthIn(nOut1_53), .SouthIn(nOut1_55), .EastIn(nOut2_54), .WestIn(nOut0_54), .ScanIn(nScanOut119), .ScanOut(nScanOut118), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_55), .NorthIn(nOut1_54), .SouthIn(nOut1_56), .EastIn(nOut2_55), .WestIn(nOut0_55), .ScanIn(nScanOut120), .ScanOut(nScanOut119), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_56), .NorthIn(nOut1_55), .SouthIn(nOut1_57), .EastIn(nOut2_56), .WestIn(nOut0_56), .ScanIn(nScanOut121), .ScanOut(nScanOut120), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_57), .NorthIn(nOut1_56), .SouthIn(nOut1_58), .EastIn(nOut2_57), .WestIn(nOut0_57), .ScanIn(nScanOut122), .ScanOut(nScanOut121), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_58), .NorthIn(nOut1_57), .SouthIn(nOut1_59), .EastIn(nOut2_58), .WestIn(nOut0_58), .ScanIn(nScanOut123), .ScanOut(nScanOut122), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_59), .NorthIn(nOut1_58), .SouthIn(nOut1_60), .EastIn(nOut2_59), .WestIn(nOut0_59), .ScanIn(nScanOut124), .ScanOut(nScanOut123), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_60), .NorthIn(nOut1_59), .SouthIn(nOut1_61), .EastIn(nOut2_60), .WestIn(nOut0_60), .ScanIn(nScanOut125), .ScanOut(nScanOut124), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_61), .NorthIn(nOut1_60), .SouthIn(nOut1_62), .EastIn(nOut2_61), .WestIn(nOut0_61), .ScanIn(nScanOut126), .ScanOut(nScanOut125), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_62), .NorthIn(nOut1_61), .SouthIn(nOut1_63), .EastIn(nOut2_62), .WestIn(nOut0_62), .ScanIn(nScanOut127), .ScanOut(nScanOut126), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_63), .ScanIn(nScanOut128), .ScanOut(nScanOut127), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_0), .ScanIn(nScanOut129), .ScanOut(nScanOut128), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_1), .NorthIn(nOut2_0), .SouthIn(nOut2_2), .EastIn(nOut3_1), .WestIn(nOut1_1), .ScanIn(nScanOut130), .ScanOut(nScanOut129), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_2), .NorthIn(nOut2_1), .SouthIn(nOut2_3), .EastIn(nOut3_2), .WestIn(nOut1_2), .ScanIn(nScanOut131), .ScanOut(nScanOut130), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_3), .NorthIn(nOut2_2), .SouthIn(nOut2_4), .EastIn(nOut3_3), .WestIn(nOut1_3), .ScanIn(nScanOut132), .ScanOut(nScanOut131), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_4), .NorthIn(nOut2_3), .SouthIn(nOut2_5), .EastIn(nOut3_4), .WestIn(nOut1_4), .ScanIn(nScanOut133), .ScanOut(nScanOut132), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_5), .NorthIn(nOut2_4), .SouthIn(nOut2_6), .EastIn(nOut3_5), .WestIn(nOut1_5), .ScanIn(nScanOut134), .ScanOut(nScanOut133), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_6), .NorthIn(nOut2_5), .SouthIn(nOut2_7), .EastIn(nOut3_6), .WestIn(nOut1_6), .ScanIn(nScanOut135), .ScanOut(nScanOut134), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_7), .NorthIn(nOut2_6), .SouthIn(nOut2_8), .EastIn(nOut3_7), .WestIn(nOut1_7), .ScanIn(nScanOut136), .ScanOut(nScanOut135), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_8), .NorthIn(nOut2_7), .SouthIn(nOut2_9), .EastIn(nOut3_8), .WestIn(nOut1_8), .ScanIn(nScanOut137), .ScanOut(nScanOut136), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_9), .NorthIn(nOut2_8), .SouthIn(nOut2_10), .EastIn(nOut3_9), .WestIn(nOut1_9), .ScanIn(nScanOut138), .ScanOut(nScanOut137), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_10), .NorthIn(nOut2_9), .SouthIn(nOut2_11), .EastIn(nOut3_10), .WestIn(nOut1_10), .ScanIn(nScanOut139), .ScanOut(nScanOut138), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_11), .NorthIn(nOut2_10), .SouthIn(nOut2_12), .EastIn(nOut3_11), .WestIn(nOut1_11), .ScanIn(nScanOut140), .ScanOut(nScanOut139), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_12), .NorthIn(nOut2_11), .SouthIn(nOut2_13), .EastIn(nOut3_12), .WestIn(nOut1_12), .ScanIn(nScanOut141), .ScanOut(nScanOut140), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_13), .NorthIn(nOut2_12), .SouthIn(nOut2_14), .EastIn(nOut3_13), .WestIn(nOut1_13), .ScanIn(nScanOut142), .ScanOut(nScanOut141), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_14), .NorthIn(nOut2_13), .SouthIn(nOut2_15), .EastIn(nOut3_14), .WestIn(nOut1_14), .ScanIn(nScanOut143), .ScanOut(nScanOut142), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_15), .NorthIn(nOut2_14), .SouthIn(nOut2_16), .EastIn(nOut3_15), .WestIn(nOut1_15), .ScanIn(nScanOut144), .ScanOut(nScanOut143), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_16), .NorthIn(nOut2_15), .SouthIn(nOut2_17), .EastIn(nOut3_16), .WestIn(nOut1_16), .ScanIn(nScanOut145), .ScanOut(nScanOut144), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_17), .NorthIn(nOut2_16), .SouthIn(nOut2_18), .EastIn(nOut3_17), .WestIn(nOut1_17), .ScanIn(nScanOut146), .ScanOut(nScanOut145), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_18), .NorthIn(nOut2_17), .SouthIn(nOut2_19), .EastIn(nOut3_18), .WestIn(nOut1_18), .ScanIn(nScanOut147), .ScanOut(nScanOut146), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_19), .NorthIn(nOut2_18), .SouthIn(nOut2_20), .EastIn(nOut3_19), .WestIn(nOut1_19), .ScanIn(nScanOut148), .ScanOut(nScanOut147), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_20), .NorthIn(nOut2_19), .SouthIn(nOut2_21), .EastIn(nOut3_20), .WestIn(nOut1_20), .ScanIn(nScanOut149), .ScanOut(nScanOut148), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_21), .NorthIn(nOut2_20), .SouthIn(nOut2_22), .EastIn(nOut3_21), .WestIn(nOut1_21), .ScanIn(nScanOut150), .ScanOut(nScanOut149), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_22), .NorthIn(nOut2_21), .SouthIn(nOut2_23), .EastIn(nOut3_22), .WestIn(nOut1_22), .ScanIn(nScanOut151), .ScanOut(nScanOut150), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_23), .NorthIn(nOut2_22), .SouthIn(nOut2_24), .EastIn(nOut3_23), .WestIn(nOut1_23), .ScanIn(nScanOut152), .ScanOut(nScanOut151), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_24), .NorthIn(nOut2_23), .SouthIn(nOut2_25), .EastIn(nOut3_24), .WestIn(nOut1_24), .ScanIn(nScanOut153), .ScanOut(nScanOut152), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_25), .NorthIn(nOut2_24), .SouthIn(nOut2_26), .EastIn(nOut3_25), .WestIn(nOut1_25), .ScanIn(nScanOut154), .ScanOut(nScanOut153), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_26), .NorthIn(nOut2_25), .SouthIn(nOut2_27), .EastIn(nOut3_26), .WestIn(nOut1_26), .ScanIn(nScanOut155), .ScanOut(nScanOut154), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_27), .NorthIn(nOut2_26), .SouthIn(nOut2_28), .EastIn(nOut3_27), .WestIn(nOut1_27), .ScanIn(nScanOut156), .ScanOut(nScanOut155), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_28), .NorthIn(nOut2_27), .SouthIn(nOut2_29), .EastIn(nOut3_28), .WestIn(nOut1_28), .ScanIn(nScanOut157), .ScanOut(nScanOut156), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_29), .NorthIn(nOut2_28), .SouthIn(nOut2_30), .EastIn(nOut3_29), .WestIn(nOut1_29), .ScanIn(nScanOut158), .ScanOut(nScanOut157), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_30), .NorthIn(nOut2_29), .SouthIn(nOut2_31), .EastIn(nOut3_30), .WestIn(nOut1_30), .ScanIn(nScanOut159), .ScanOut(nScanOut158), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_31), .NorthIn(nOut2_30), .SouthIn(nOut2_32), .EastIn(nOut3_31), .WestIn(nOut1_31), .ScanIn(nScanOut160), .ScanOut(nScanOut159), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_32), .NorthIn(nOut2_31), .SouthIn(nOut2_33), .EastIn(nOut3_32), .WestIn(nOut1_32), .ScanIn(nScanOut161), .ScanOut(nScanOut160), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_33), .NorthIn(nOut2_32), .SouthIn(nOut2_34), .EastIn(nOut3_33), .WestIn(nOut1_33), .ScanIn(nScanOut162), .ScanOut(nScanOut161), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_34), .NorthIn(nOut2_33), .SouthIn(nOut2_35), .EastIn(nOut3_34), .WestIn(nOut1_34), .ScanIn(nScanOut163), .ScanOut(nScanOut162), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_35), .NorthIn(nOut2_34), .SouthIn(nOut2_36), .EastIn(nOut3_35), .WestIn(nOut1_35), .ScanIn(nScanOut164), .ScanOut(nScanOut163), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_36), .NorthIn(nOut2_35), .SouthIn(nOut2_37), .EastIn(nOut3_36), .WestIn(nOut1_36), .ScanIn(nScanOut165), .ScanOut(nScanOut164), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_37), .NorthIn(nOut2_36), .SouthIn(nOut2_38), .EastIn(nOut3_37), .WestIn(nOut1_37), .ScanIn(nScanOut166), .ScanOut(nScanOut165), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_38), .NorthIn(nOut2_37), .SouthIn(nOut2_39), .EastIn(nOut3_38), .WestIn(nOut1_38), .ScanIn(nScanOut167), .ScanOut(nScanOut166), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_39), .NorthIn(nOut2_38), .SouthIn(nOut2_40), .EastIn(nOut3_39), .WestIn(nOut1_39), .ScanIn(nScanOut168), .ScanOut(nScanOut167), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_40), .NorthIn(nOut2_39), .SouthIn(nOut2_41), .EastIn(nOut3_40), .WestIn(nOut1_40), .ScanIn(nScanOut169), .ScanOut(nScanOut168), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_41), .NorthIn(nOut2_40), .SouthIn(nOut2_42), .EastIn(nOut3_41), .WestIn(nOut1_41), .ScanIn(nScanOut170), .ScanOut(nScanOut169), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_42), .NorthIn(nOut2_41), .SouthIn(nOut2_43), .EastIn(nOut3_42), .WestIn(nOut1_42), .ScanIn(nScanOut171), .ScanOut(nScanOut170), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_43), .NorthIn(nOut2_42), .SouthIn(nOut2_44), .EastIn(nOut3_43), .WestIn(nOut1_43), .ScanIn(nScanOut172), .ScanOut(nScanOut171), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_44), .NorthIn(nOut2_43), .SouthIn(nOut2_45), .EastIn(nOut3_44), .WestIn(nOut1_44), .ScanIn(nScanOut173), .ScanOut(nScanOut172), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_45), .NorthIn(nOut2_44), .SouthIn(nOut2_46), .EastIn(nOut3_45), .WestIn(nOut1_45), .ScanIn(nScanOut174), .ScanOut(nScanOut173), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_46), .NorthIn(nOut2_45), .SouthIn(nOut2_47), .EastIn(nOut3_46), .WestIn(nOut1_46), .ScanIn(nScanOut175), .ScanOut(nScanOut174), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_47), .NorthIn(nOut2_46), .SouthIn(nOut2_48), .EastIn(nOut3_47), .WestIn(nOut1_47), .ScanIn(nScanOut176), .ScanOut(nScanOut175), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_48), .NorthIn(nOut2_47), .SouthIn(nOut2_49), .EastIn(nOut3_48), .WestIn(nOut1_48), .ScanIn(nScanOut177), .ScanOut(nScanOut176), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_49), .NorthIn(nOut2_48), .SouthIn(nOut2_50), .EastIn(nOut3_49), .WestIn(nOut1_49), .ScanIn(nScanOut178), .ScanOut(nScanOut177), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_50), .NorthIn(nOut2_49), .SouthIn(nOut2_51), .EastIn(nOut3_50), .WestIn(nOut1_50), .ScanIn(nScanOut179), .ScanOut(nScanOut178), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_51), .NorthIn(nOut2_50), .SouthIn(nOut2_52), .EastIn(nOut3_51), .WestIn(nOut1_51), .ScanIn(nScanOut180), .ScanOut(nScanOut179), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_52), .NorthIn(nOut2_51), .SouthIn(nOut2_53), .EastIn(nOut3_52), .WestIn(nOut1_52), .ScanIn(nScanOut181), .ScanOut(nScanOut180), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_53), .NorthIn(nOut2_52), .SouthIn(nOut2_54), .EastIn(nOut3_53), .WestIn(nOut1_53), .ScanIn(nScanOut182), .ScanOut(nScanOut181), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_54), .NorthIn(nOut2_53), .SouthIn(nOut2_55), .EastIn(nOut3_54), .WestIn(nOut1_54), .ScanIn(nScanOut183), .ScanOut(nScanOut182), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_55), .NorthIn(nOut2_54), .SouthIn(nOut2_56), .EastIn(nOut3_55), .WestIn(nOut1_55), .ScanIn(nScanOut184), .ScanOut(nScanOut183), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_56), .NorthIn(nOut2_55), .SouthIn(nOut2_57), .EastIn(nOut3_56), .WestIn(nOut1_56), .ScanIn(nScanOut185), .ScanOut(nScanOut184), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_57), .NorthIn(nOut2_56), .SouthIn(nOut2_58), .EastIn(nOut3_57), .WestIn(nOut1_57), .ScanIn(nScanOut186), .ScanOut(nScanOut185), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_58), .NorthIn(nOut2_57), .SouthIn(nOut2_59), .EastIn(nOut3_58), .WestIn(nOut1_58), .ScanIn(nScanOut187), .ScanOut(nScanOut186), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_59), .NorthIn(nOut2_58), .SouthIn(nOut2_60), .EastIn(nOut3_59), .WestIn(nOut1_59), .ScanIn(nScanOut188), .ScanOut(nScanOut187), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_60), .NorthIn(nOut2_59), .SouthIn(nOut2_61), .EastIn(nOut3_60), .WestIn(nOut1_60), .ScanIn(nScanOut189), .ScanOut(nScanOut188), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_61), .NorthIn(nOut2_60), .SouthIn(nOut2_62), .EastIn(nOut3_61), .WestIn(nOut1_61), .ScanIn(nScanOut190), .ScanOut(nScanOut189), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_62), .NorthIn(nOut2_61), .SouthIn(nOut2_63), .EastIn(nOut3_62), .WestIn(nOut1_62), .ScanIn(nScanOut191), .ScanOut(nScanOut190), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_63), .ScanIn(nScanOut192), .ScanOut(nScanOut191), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_0), .ScanIn(nScanOut193), .ScanOut(nScanOut192), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_1), .NorthIn(nOut3_0), .SouthIn(nOut3_2), .EastIn(nOut4_1), .WestIn(nOut2_1), .ScanIn(nScanOut194), .ScanOut(nScanOut193), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_2), .NorthIn(nOut3_1), .SouthIn(nOut3_3), .EastIn(nOut4_2), .WestIn(nOut2_2), .ScanIn(nScanOut195), .ScanOut(nScanOut194), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_3), .NorthIn(nOut3_2), .SouthIn(nOut3_4), .EastIn(nOut4_3), .WestIn(nOut2_3), .ScanIn(nScanOut196), .ScanOut(nScanOut195), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_4), .NorthIn(nOut3_3), .SouthIn(nOut3_5), .EastIn(nOut4_4), .WestIn(nOut2_4), .ScanIn(nScanOut197), .ScanOut(nScanOut196), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_5), .NorthIn(nOut3_4), .SouthIn(nOut3_6), .EastIn(nOut4_5), .WestIn(nOut2_5), .ScanIn(nScanOut198), .ScanOut(nScanOut197), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_6), .NorthIn(nOut3_5), .SouthIn(nOut3_7), .EastIn(nOut4_6), .WestIn(nOut2_6), .ScanIn(nScanOut199), .ScanOut(nScanOut198), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_7), .NorthIn(nOut3_6), .SouthIn(nOut3_8), .EastIn(nOut4_7), .WestIn(nOut2_7), .ScanIn(nScanOut200), .ScanOut(nScanOut199), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_8), .NorthIn(nOut3_7), .SouthIn(nOut3_9), .EastIn(nOut4_8), .WestIn(nOut2_8), .ScanIn(nScanOut201), .ScanOut(nScanOut200), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_9), .NorthIn(nOut3_8), .SouthIn(nOut3_10), .EastIn(nOut4_9), .WestIn(nOut2_9), .ScanIn(nScanOut202), .ScanOut(nScanOut201), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_10), .NorthIn(nOut3_9), .SouthIn(nOut3_11), .EastIn(nOut4_10), .WestIn(nOut2_10), .ScanIn(nScanOut203), .ScanOut(nScanOut202), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_11), .NorthIn(nOut3_10), .SouthIn(nOut3_12), .EastIn(nOut4_11), .WestIn(nOut2_11), .ScanIn(nScanOut204), .ScanOut(nScanOut203), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_12), .NorthIn(nOut3_11), .SouthIn(nOut3_13), .EastIn(nOut4_12), .WestIn(nOut2_12), .ScanIn(nScanOut205), .ScanOut(nScanOut204), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_13), .NorthIn(nOut3_12), .SouthIn(nOut3_14), .EastIn(nOut4_13), .WestIn(nOut2_13), .ScanIn(nScanOut206), .ScanOut(nScanOut205), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_14), .NorthIn(nOut3_13), .SouthIn(nOut3_15), .EastIn(nOut4_14), .WestIn(nOut2_14), .ScanIn(nScanOut207), .ScanOut(nScanOut206), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_15), .NorthIn(nOut3_14), .SouthIn(nOut3_16), .EastIn(nOut4_15), .WestIn(nOut2_15), .ScanIn(nScanOut208), .ScanOut(nScanOut207), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_16), .NorthIn(nOut3_15), .SouthIn(nOut3_17), .EastIn(nOut4_16), .WestIn(nOut2_16), .ScanIn(nScanOut209), .ScanOut(nScanOut208), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_17), .NorthIn(nOut3_16), .SouthIn(nOut3_18), .EastIn(nOut4_17), .WestIn(nOut2_17), .ScanIn(nScanOut210), .ScanOut(nScanOut209), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_18), .NorthIn(nOut3_17), .SouthIn(nOut3_19), .EastIn(nOut4_18), .WestIn(nOut2_18), .ScanIn(nScanOut211), .ScanOut(nScanOut210), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_19), .NorthIn(nOut3_18), .SouthIn(nOut3_20), .EastIn(nOut4_19), .WestIn(nOut2_19), .ScanIn(nScanOut212), .ScanOut(nScanOut211), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_20), .NorthIn(nOut3_19), .SouthIn(nOut3_21), .EastIn(nOut4_20), .WestIn(nOut2_20), .ScanIn(nScanOut213), .ScanOut(nScanOut212), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_21), .NorthIn(nOut3_20), .SouthIn(nOut3_22), .EastIn(nOut4_21), .WestIn(nOut2_21), .ScanIn(nScanOut214), .ScanOut(nScanOut213), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_22), .NorthIn(nOut3_21), .SouthIn(nOut3_23), .EastIn(nOut4_22), .WestIn(nOut2_22), .ScanIn(nScanOut215), .ScanOut(nScanOut214), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_23), .NorthIn(nOut3_22), .SouthIn(nOut3_24), .EastIn(nOut4_23), .WestIn(nOut2_23), .ScanIn(nScanOut216), .ScanOut(nScanOut215), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_24), .NorthIn(nOut3_23), .SouthIn(nOut3_25), .EastIn(nOut4_24), .WestIn(nOut2_24), .ScanIn(nScanOut217), .ScanOut(nScanOut216), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_25), .NorthIn(nOut3_24), .SouthIn(nOut3_26), .EastIn(nOut4_25), .WestIn(nOut2_25), .ScanIn(nScanOut218), .ScanOut(nScanOut217), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_26), .NorthIn(nOut3_25), .SouthIn(nOut3_27), .EastIn(nOut4_26), .WestIn(nOut2_26), .ScanIn(nScanOut219), .ScanOut(nScanOut218), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_27), .NorthIn(nOut3_26), .SouthIn(nOut3_28), .EastIn(nOut4_27), .WestIn(nOut2_27), .ScanIn(nScanOut220), .ScanOut(nScanOut219), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_28), .NorthIn(nOut3_27), .SouthIn(nOut3_29), .EastIn(nOut4_28), .WestIn(nOut2_28), .ScanIn(nScanOut221), .ScanOut(nScanOut220), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_29), .NorthIn(nOut3_28), .SouthIn(nOut3_30), .EastIn(nOut4_29), .WestIn(nOut2_29), .ScanIn(nScanOut222), .ScanOut(nScanOut221), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_30), .NorthIn(nOut3_29), .SouthIn(nOut3_31), .EastIn(nOut4_30), .WestIn(nOut2_30), .ScanIn(nScanOut223), .ScanOut(nScanOut222), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_31), .NorthIn(nOut3_30), .SouthIn(nOut3_32), .EastIn(nOut4_31), .WestIn(nOut2_31), .ScanIn(nScanOut224), .ScanOut(nScanOut223), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_32), .NorthIn(nOut3_31), .SouthIn(nOut3_33), .EastIn(nOut4_32), .WestIn(nOut2_32), .ScanIn(nScanOut225), .ScanOut(nScanOut224), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_33), .NorthIn(nOut3_32), .SouthIn(nOut3_34), .EastIn(nOut4_33), .WestIn(nOut2_33), .ScanIn(nScanOut226), .ScanOut(nScanOut225), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_34), .NorthIn(nOut3_33), .SouthIn(nOut3_35), .EastIn(nOut4_34), .WestIn(nOut2_34), .ScanIn(nScanOut227), .ScanOut(nScanOut226), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_35), .NorthIn(nOut3_34), .SouthIn(nOut3_36), .EastIn(nOut4_35), .WestIn(nOut2_35), .ScanIn(nScanOut228), .ScanOut(nScanOut227), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_36), .NorthIn(nOut3_35), .SouthIn(nOut3_37), .EastIn(nOut4_36), .WestIn(nOut2_36), .ScanIn(nScanOut229), .ScanOut(nScanOut228), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_37), .NorthIn(nOut3_36), .SouthIn(nOut3_38), .EastIn(nOut4_37), .WestIn(nOut2_37), .ScanIn(nScanOut230), .ScanOut(nScanOut229), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_38), .NorthIn(nOut3_37), .SouthIn(nOut3_39), .EastIn(nOut4_38), .WestIn(nOut2_38), .ScanIn(nScanOut231), .ScanOut(nScanOut230), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_39), .NorthIn(nOut3_38), .SouthIn(nOut3_40), .EastIn(nOut4_39), .WestIn(nOut2_39), .ScanIn(nScanOut232), .ScanOut(nScanOut231), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_40), .NorthIn(nOut3_39), .SouthIn(nOut3_41), .EastIn(nOut4_40), .WestIn(nOut2_40), .ScanIn(nScanOut233), .ScanOut(nScanOut232), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_41), .NorthIn(nOut3_40), .SouthIn(nOut3_42), .EastIn(nOut4_41), .WestIn(nOut2_41), .ScanIn(nScanOut234), .ScanOut(nScanOut233), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_42), .NorthIn(nOut3_41), .SouthIn(nOut3_43), .EastIn(nOut4_42), .WestIn(nOut2_42), .ScanIn(nScanOut235), .ScanOut(nScanOut234), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_43), .NorthIn(nOut3_42), .SouthIn(nOut3_44), .EastIn(nOut4_43), .WestIn(nOut2_43), .ScanIn(nScanOut236), .ScanOut(nScanOut235), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_44), .NorthIn(nOut3_43), .SouthIn(nOut3_45), .EastIn(nOut4_44), .WestIn(nOut2_44), .ScanIn(nScanOut237), .ScanOut(nScanOut236), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_45), .NorthIn(nOut3_44), .SouthIn(nOut3_46), .EastIn(nOut4_45), .WestIn(nOut2_45), .ScanIn(nScanOut238), .ScanOut(nScanOut237), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_46), .NorthIn(nOut3_45), .SouthIn(nOut3_47), .EastIn(nOut4_46), .WestIn(nOut2_46), .ScanIn(nScanOut239), .ScanOut(nScanOut238), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_47), .NorthIn(nOut3_46), .SouthIn(nOut3_48), .EastIn(nOut4_47), .WestIn(nOut2_47), .ScanIn(nScanOut240), .ScanOut(nScanOut239), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_48), .NorthIn(nOut3_47), .SouthIn(nOut3_49), .EastIn(nOut4_48), .WestIn(nOut2_48), .ScanIn(nScanOut241), .ScanOut(nScanOut240), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_49), .NorthIn(nOut3_48), .SouthIn(nOut3_50), .EastIn(nOut4_49), .WestIn(nOut2_49), .ScanIn(nScanOut242), .ScanOut(nScanOut241), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_50), .NorthIn(nOut3_49), .SouthIn(nOut3_51), .EastIn(nOut4_50), .WestIn(nOut2_50), .ScanIn(nScanOut243), .ScanOut(nScanOut242), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_51), .NorthIn(nOut3_50), .SouthIn(nOut3_52), .EastIn(nOut4_51), .WestIn(nOut2_51), .ScanIn(nScanOut244), .ScanOut(nScanOut243), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_52), .NorthIn(nOut3_51), .SouthIn(nOut3_53), .EastIn(nOut4_52), .WestIn(nOut2_52), .ScanIn(nScanOut245), .ScanOut(nScanOut244), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_53), .NorthIn(nOut3_52), .SouthIn(nOut3_54), .EastIn(nOut4_53), .WestIn(nOut2_53), .ScanIn(nScanOut246), .ScanOut(nScanOut245), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_54), .NorthIn(nOut3_53), .SouthIn(nOut3_55), .EastIn(nOut4_54), .WestIn(nOut2_54), .ScanIn(nScanOut247), .ScanOut(nScanOut246), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_55), .NorthIn(nOut3_54), .SouthIn(nOut3_56), .EastIn(nOut4_55), .WestIn(nOut2_55), .ScanIn(nScanOut248), .ScanOut(nScanOut247), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_56), .NorthIn(nOut3_55), .SouthIn(nOut3_57), .EastIn(nOut4_56), .WestIn(nOut2_56), .ScanIn(nScanOut249), .ScanOut(nScanOut248), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_57), .NorthIn(nOut3_56), .SouthIn(nOut3_58), .EastIn(nOut4_57), .WestIn(nOut2_57), .ScanIn(nScanOut250), .ScanOut(nScanOut249), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_58), .NorthIn(nOut3_57), .SouthIn(nOut3_59), .EastIn(nOut4_58), .WestIn(nOut2_58), .ScanIn(nScanOut251), .ScanOut(nScanOut250), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_59), .NorthIn(nOut3_58), .SouthIn(nOut3_60), .EastIn(nOut4_59), .WestIn(nOut2_59), .ScanIn(nScanOut252), .ScanOut(nScanOut251), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_60), .NorthIn(nOut3_59), .SouthIn(nOut3_61), .EastIn(nOut4_60), .WestIn(nOut2_60), .ScanIn(nScanOut253), .ScanOut(nScanOut252), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_61), .NorthIn(nOut3_60), .SouthIn(nOut3_62), .EastIn(nOut4_61), .WestIn(nOut2_61), .ScanIn(nScanOut254), .ScanOut(nScanOut253), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_62), .NorthIn(nOut3_61), .SouthIn(nOut3_63), .EastIn(nOut4_62), .WestIn(nOut2_62), .ScanIn(nScanOut255), .ScanOut(nScanOut254), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_63), .ScanIn(nScanOut256), .ScanOut(nScanOut255), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_256 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_0), .ScanIn(nScanOut257), .ScanOut(nScanOut256), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_257 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_1), .NorthIn(nOut4_0), .SouthIn(nOut4_2), .EastIn(nOut5_1), .WestIn(nOut3_1), .ScanIn(nScanOut258), .ScanOut(nScanOut257), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_258 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_2), .NorthIn(nOut4_1), .SouthIn(nOut4_3), .EastIn(nOut5_2), .WestIn(nOut3_2), .ScanIn(nScanOut259), .ScanOut(nScanOut258), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_259 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_3), .NorthIn(nOut4_2), .SouthIn(nOut4_4), .EastIn(nOut5_3), .WestIn(nOut3_3), .ScanIn(nScanOut260), .ScanOut(nScanOut259), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_260 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_4), .NorthIn(nOut4_3), .SouthIn(nOut4_5), .EastIn(nOut5_4), .WestIn(nOut3_4), .ScanIn(nScanOut261), .ScanOut(nScanOut260), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_261 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_5), .NorthIn(nOut4_4), .SouthIn(nOut4_6), .EastIn(nOut5_5), .WestIn(nOut3_5), .ScanIn(nScanOut262), .ScanOut(nScanOut261), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_262 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_6), .NorthIn(nOut4_5), .SouthIn(nOut4_7), .EastIn(nOut5_6), .WestIn(nOut3_6), .ScanIn(nScanOut263), .ScanOut(nScanOut262), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_263 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_7), .NorthIn(nOut4_6), .SouthIn(nOut4_8), .EastIn(nOut5_7), .WestIn(nOut3_7), .ScanIn(nScanOut264), .ScanOut(nScanOut263), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_264 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_8), .NorthIn(nOut4_7), .SouthIn(nOut4_9), .EastIn(nOut5_8), .WestIn(nOut3_8), .ScanIn(nScanOut265), .ScanOut(nScanOut264), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_265 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_9), .NorthIn(nOut4_8), .SouthIn(nOut4_10), .EastIn(nOut5_9), .WestIn(nOut3_9), .ScanIn(nScanOut266), .ScanOut(nScanOut265), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_266 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_10), .NorthIn(nOut4_9), .SouthIn(nOut4_11), .EastIn(nOut5_10), .WestIn(nOut3_10), .ScanIn(nScanOut267), .ScanOut(nScanOut266), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_267 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_11), .NorthIn(nOut4_10), .SouthIn(nOut4_12), .EastIn(nOut5_11), .WestIn(nOut3_11), .ScanIn(nScanOut268), .ScanOut(nScanOut267), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_268 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_12), .NorthIn(nOut4_11), .SouthIn(nOut4_13), .EastIn(nOut5_12), .WestIn(nOut3_12), .ScanIn(nScanOut269), .ScanOut(nScanOut268), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_269 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_13), .NorthIn(nOut4_12), .SouthIn(nOut4_14), .EastIn(nOut5_13), .WestIn(nOut3_13), .ScanIn(nScanOut270), .ScanOut(nScanOut269), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_270 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_14), .NorthIn(nOut4_13), .SouthIn(nOut4_15), .EastIn(nOut5_14), .WestIn(nOut3_14), .ScanIn(nScanOut271), .ScanOut(nScanOut270), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_271 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_15), .NorthIn(nOut4_14), .SouthIn(nOut4_16), .EastIn(nOut5_15), .WestIn(nOut3_15), .ScanIn(nScanOut272), .ScanOut(nScanOut271), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_272 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_16), .NorthIn(nOut4_15), .SouthIn(nOut4_17), .EastIn(nOut5_16), .WestIn(nOut3_16), .ScanIn(nScanOut273), .ScanOut(nScanOut272), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_273 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_17), .NorthIn(nOut4_16), .SouthIn(nOut4_18), .EastIn(nOut5_17), .WestIn(nOut3_17), .ScanIn(nScanOut274), .ScanOut(nScanOut273), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_274 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_18), .NorthIn(nOut4_17), .SouthIn(nOut4_19), .EastIn(nOut5_18), .WestIn(nOut3_18), .ScanIn(nScanOut275), .ScanOut(nScanOut274), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_275 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_19), .NorthIn(nOut4_18), .SouthIn(nOut4_20), .EastIn(nOut5_19), .WestIn(nOut3_19), .ScanIn(nScanOut276), .ScanOut(nScanOut275), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_276 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_20), .NorthIn(nOut4_19), .SouthIn(nOut4_21), .EastIn(nOut5_20), .WestIn(nOut3_20), .ScanIn(nScanOut277), .ScanOut(nScanOut276), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_277 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_21), .NorthIn(nOut4_20), .SouthIn(nOut4_22), .EastIn(nOut5_21), .WestIn(nOut3_21), .ScanIn(nScanOut278), .ScanOut(nScanOut277), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_278 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_22), .NorthIn(nOut4_21), .SouthIn(nOut4_23), .EastIn(nOut5_22), .WestIn(nOut3_22), .ScanIn(nScanOut279), .ScanOut(nScanOut278), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_279 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_23), .NorthIn(nOut4_22), .SouthIn(nOut4_24), .EastIn(nOut5_23), .WestIn(nOut3_23), .ScanIn(nScanOut280), .ScanOut(nScanOut279), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_280 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_24), .NorthIn(nOut4_23), .SouthIn(nOut4_25), .EastIn(nOut5_24), .WestIn(nOut3_24), .ScanIn(nScanOut281), .ScanOut(nScanOut280), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_281 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_25), .NorthIn(nOut4_24), .SouthIn(nOut4_26), .EastIn(nOut5_25), .WestIn(nOut3_25), .ScanIn(nScanOut282), .ScanOut(nScanOut281), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_282 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_26), .NorthIn(nOut4_25), .SouthIn(nOut4_27), .EastIn(nOut5_26), .WestIn(nOut3_26), .ScanIn(nScanOut283), .ScanOut(nScanOut282), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_283 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_27), .NorthIn(nOut4_26), .SouthIn(nOut4_28), .EastIn(nOut5_27), .WestIn(nOut3_27), .ScanIn(nScanOut284), .ScanOut(nScanOut283), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_284 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_28), .NorthIn(nOut4_27), .SouthIn(nOut4_29), .EastIn(nOut5_28), .WestIn(nOut3_28), .ScanIn(nScanOut285), .ScanOut(nScanOut284), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_285 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_29), .NorthIn(nOut4_28), .SouthIn(nOut4_30), .EastIn(nOut5_29), .WestIn(nOut3_29), .ScanIn(nScanOut286), .ScanOut(nScanOut285), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_286 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_30), .NorthIn(nOut4_29), .SouthIn(nOut4_31), .EastIn(nOut5_30), .WestIn(nOut3_30), .ScanIn(nScanOut287), .ScanOut(nScanOut286), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_287 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_31), .NorthIn(nOut4_30), .SouthIn(nOut4_32), .EastIn(nOut5_31), .WestIn(nOut3_31), .ScanIn(nScanOut288), .ScanOut(nScanOut287), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_288 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_32), .NorthIn(nOut4_31), .SouthIn(nOut4_33), .EastIn(nOut5_32), .WestIn(nOut3_32), .ScanIn(nScanOut289), .ScanOut(nScanOut288), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_289 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_33), .NorthIn(nOut4_32), .SouthIn(nOut4_34), .EastIn(nOut5_33), .WestIn(nOut3_33), .ScanIn(nScanOut290), .ScanOut(nScanOut289), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_290 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_34), .NorthIn(nOut4_33), .SouthIn(nOut4_35), .EastIn(nOut5_34), .WestIn(nOut3_34), .ScanIn(nScanOut291), .ScanOut(nScanOut290), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_291 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_35), .NorthIn(nOut4_34), .SouthIn(nOut4_36), .EastIn(nOut5_35), .WestIn(nOut3_35), .ScanIn(nScanOut292), .ScanOut(nScanOut291), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_292 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_36), .NorthIn(nOut4_35), .SouthIn(nOut4_37), .EastIn(nOut5_36), .WestIn(nOut3_36), .ScanIn(nScanOut293), .ScanOut(nScanOut292), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_293 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_37), .NorthIn(nOut4_36), .SouthIn(nOut4_38), .EastIn(nOut5_37), .WestIn(nOut3_37), .ScanIn(nScanOut294), .ScanOut(nScanOut293), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_294 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_38), .NorthIn(nOut4_37), .SouthIn(nOut4_39), .EastIn(nOut5_38), .WestIn(nOut3_38), .ScanIn(nScanOut295), .ScanOut(nScanOut294), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_295 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_39), .NorthIn(nOut4_38), .SouthIn(nOut4_40), .EastIn(nOut5_39), .WestIn(nOut3_39), .ScanIn(nScanOut296), .ScanOut(nScanOut295), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_296 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_40), .NorthIn(nOut4_39), .SouthIn(nOut4_41), .EastIn(nOut5_40), .WestIn(nOut3_40), .ScanIn(nScanOut297), .ScanOut(nScanOut296), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_297 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_41), .NorthIn(nOut4_40), .SouthIn(nOut4_42), .EastIn(nOut5_41), .WestIn(nOut3_41), .ScanIn(nScanOut298), .ScanOut(nScanOut297), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_298 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_42), .NorthIn(nOut4_41), .SouthIn(nOut4_43), .EastIn(nOut5_42), .WestIn(nOut3_42), .ScanIn(nScanOut299), .ScanOut(nScanOut298), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_299 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_43), .NorthIn(nOut4_42), .SouthIn(nOut4_44), .EastIn(nOut5_43), .WestIn(nOut3_43), .ScanIn(nScanOut300), .ScanOut(nScanOut299), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_300 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_44), .NorthIn(nOut4_43), .SouthIn(nOut4_45), .EastIn(nOut5_44), .WestIn(nOut3_44), .ScanIn(nScanOut301), .ScanOut(nScanOut300), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_301 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_45), .NorthIn(nOut4_44), .SouthIn(nOut4_46), .EastIn(nOut5_45), .WestIn(nOut3_45), .ScanIn(nScanOut302), .ScanOut(nScanOut301), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_302 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_46), .NorthIn(nOut4_45), .SouthIn(nOut4_47), .EastIn(nOut5_46), .WestIn(nOut3_46), .ScanIn(nScanOut303), .ScanOut(nScanOut302), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_303 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_47), .NorthIn(nOut4_46), .SouthIn(nOut4_48), .EastIn(nOut5_47), .WestIn(nOut3_47), .ScanIn(nScanOut304), .ScanOut(nScanOut303), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_304 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_48), .NorthIn(nOut4_47), .SouthIn(nOut4_49), .EastIn(nOut5_48), .WestIn(nOut3_48), .ScanIn(nScanOut305), .ScanOut(nScanOut304), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_305 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_49), .NorthIn(nOut4_48), .SouthIn(nOut4_50), .EastIn(nOut5_49), .WestIn(nOut3_49), .ScanIn(nScanOut306), .ScanOut(nScanOut305), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_306 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_50), .NorthIn(nOut4_49), .SouthIn(nOut4_51), .EastIn(nOut5_50), .WestIn(nOut3_50), .ScanIn(nScanOut307), .ScanOut(nScanOut306), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_307 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_51), .NorthIn(nOut4_50), .SouthIn(nOut4_52), .EastIn(nOut5_51), .WestIn(nOut3_51), .ScanIn(nScanOut308), .ScanOut(nScanOut307), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_308 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_52), .NorthIn(nOut4_51), .SouthIn(nOut4_53), .EastIn(nOut5_52), .WestIn(nOut3_52), .ScanIn(nScanOut309), .ScanOut(nScanOut308), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_309 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_53), .NorthIn(nOut4_52), .SouthIn(nOut4_54), .EastIn(nOut5_53), .WestIn(nOut3_53), .ScanIn(nScanOut310), .ScanOut(nScanOut309), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_310 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_54), .NorthIn(nOut4_53), .SouthIn(nOut4_55), .EastIn(nOut5_54), .WestIn(nOut3_54), .ScanIn(nScanOut311), .ScanOut(nScanOut310), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_311 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_55), .NorthIn(nOut4_54), .SouthIn(nOut4_56), .EastIn(nOut5_55), .WestIn(nOut3_55), .ScanIn(nScanOut312), .ScanOut(nScanOut311), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_312 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_56), .NorthIn(nOut4_55), .SouthIn(nOut4_57), .EastIn(nOut5_56), .WestIn(nOut3_56), .ScanIn(nScanOut313), .ScanOut(nScanOut312), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_313 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_57), .NorthIn(nOut4_56), .SouthIn(nOut4_58), .EastIn(nOut5_57), .WestIn(nOut3_57), .ScanIn(nScanOut314), .ScanOut(nScanOut313), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_314 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_58), .NorthIn(nOut4_57), .SouthIn(nOut4_59), .EastIn(nOut5_58), .WestIn(nOut3_58), .ScanIn(nScanOut315), .ScanOut(nScanOut314), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_315 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_59), .NorthIn(nOut4_58), .SouthIn(nOut4_60), .EastIn(nOut5_59), .WestIn(nOut3_59), .ScanIn(nScanOut316), .ScanOut(nScanOut315), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_316 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_60), .NorthIn(nOut4_59), .SouthIn(nOut4_61), .EastIn(nOut5_60), .WestIn(nOut3_60), .ScanIn(nScanOut317), .ScanOut(nScanOut316), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_317 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_61), .NorthIn(nOut4_60), .SouthIn(nOut4_62), .EastIn(nOut5_61), .WestIn(nOut3_61), .ScanIn(nScanOut318), .ScanOut(nScanOut317), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_318 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_62), .NorthIn(nOut4_61), .SouthIn(nOut4_63), .EastIn(nOut5_62), .WestIn(nOut3_62), .ScanIn(nScanOut319), .ScanOut(nScanOut318), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_319 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_63), .ScanIn(nScanOut320), .ScanOut(nScanOut319), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_320 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_0), .ScanIn(nScanOut321), .ScanOut(nScanOut320), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_321 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_1), .NorthIn(nOut5_0), .SouthIn(nOut5_2), .EastIn(nOut6_1), .WestIn(nOut4_1), .ScanIn(nScanOut322), .ScanOut(nScanOut321), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_322 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_2), .NorthIn(nOut5_1), .SouthIn(nOut5_3), .EastIn(nOut6_2), .WestIn(nOut4_2), .ScanIn(nScanOut323), .ScanOut(nScanOut322), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_323 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_3), .NorthIn(nOut5_2), .SouthIn(nOut5_4), .EastIn(nOut6_3), .WestIn(nOut4_3), .ScanIn(nScanOut324), .ScanOut(nScanOut323), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_324 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_4), .NorthIn(nOut5_3), .SouthIn(nOut5_5), .EastIn(nOut6_4), .WestIn(nOut4_4), .ScanIn(nScanOut325), .ScanOut(nScanOut324), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_325 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_5), .NorthIn(nOut5_4), .SouthIn(nOut5_6), .EastIn(nOut6_5), .WestIn(nOut4_5), .ScanIn(nScanOut326), .ScanOut(nScanOut325), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_326 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_6), .NorthIn(nOut5_5), .SouthIn(nOut5_7), .EastIn(nOut6_6), .WestIn(nOut4_6), .ScanIn(nScanOut327), .ScanOut(nScanOut326), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_327 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_7), .NorthIn(nOut5_6), .SouthIn(nOut5_8), .EastIn(nOut6_7), .WestIn(nOut4_7), .ScanIn(nScanOut328), .ScanOut(nScanOut327), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_328 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_8), .NorthIn(nOut5_7), .SouthIn(nOut5_9), .EastIn(nOut6_8), .WestIn(nOut4_8), .ScanIn(nScanOut329), .ScanOut(nScanOut328), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_329 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_9), .NorthIn(nOut5_8), .SouthIn(nOut5_10), .EastIn(nOut6_9), .WestIn(nOut4_9), .ScanIn(nScanOut330), .ScanOut(nScanOut329), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_330 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_10), .NorthIn(nOut5_9), .SouthIn(nOut5_11), .EastIn(nOut6_10), .WestIn(nOut4_10), .ScanIn(nScanOut331), .ScanOut(nScanOut330), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_331 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_11), .NorthIn(nOut5_10), .SouthIn(nOut5_12), .EastIn(nOut6_11), .WestIn(nOut4_11), .ScanIn(nScanOut332), .ScanOut(nScanOut331), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_332 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_12), .NorthIn(nOut5_11), .SouthIn(nOut5_13), .EastIn(nOut6_12), .WestIn(nOut4_12), .ScanIn(nScanOut333), .ScanOut(nScanOut332), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_333 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_13), .NorthIn(nOut5_12), .SouthIn(nOut5_14), .EastIn(nOut6_13), .WestIn(nOut4_13), .ScanIn(nScanOut334), .ScanOut(nScanOut333), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_334 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_14), .NorthIn(nOut5_13), .SouthIn(nOut5_15), .EastIn(nOut6_14), .WestIn(nOut4_14), .ScanIn(nScanOut335), .ScanOut(nScanOut334), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_335 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_15), .NorthIn(nOut5_14), .SouthIn(nOut5_16), .EastIn(nOut6_15), .WestIn(nOut4_15), .ScanIn(nScanOut336), .ScanOut(nScanOut335), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_336 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_16), .NorthIn(nOut5_15), .SouthIn(nOut5_17), .EastIn(nOut6_16), .WestIn(nOut4_16), .ScanIn(nScanOut337), .ScanOut(nScanOut336), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_337 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_17), .NorthIn(nOut5_16), .SouthIn(nOut5_18), .EastIn(nOut6_17), .WestIn(nOut4_17), .ScanIn(nScanOut338), .ScanOut(nScanOut337), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_338 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_18), .NorthIn(nOut5_17), .SouthIn(nOut5_19), .EastIn(nOut6_18), .WestIn(nOut4_18), .ScanIn(nScanOut339), .ScanOut(nScanOut338), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_339 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_19), .NorthIn(nOut5_18), .SouthIn(nOut5_20), .EastIn(nOut6_19), .WestIn(nOut4_19), .ScanIn(nScanOut340), .ScanOut(nScanOut339), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_340 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_20), .NorthIn(nOut5_19), .SouthIn(nOut5_21), .EastIn(nOut6_20), .WestIn(nOut4_20), .ScanIn(nScanOut341), .ScanOut(nScanOut340), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_341 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_21), .NorthIn(nOut5_20), .SouthIn(nOut5_22), .EastIn(nOut6_21), .WestIn(nOut4_21), .ScanIn(nScanOut342), .ScanOut(nScanOut341), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_342 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_22), .NorthIn(nOut5_21), .SouthIn(nOut5_23), .EastIn(nOut6_22), .WestIn(nOut4_22), .ScanIn(nScanOut343), .ScanOut(nScanOut342), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_343 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_23), .NorthIn(nOut5_22), .SouthIn(nOut5_24), .EastIn(nOut6_23), .WestIn(nOut4_23), .ScanIn(nScanOut344), .ScanOut(nScanOut343), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_344 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_24), .NorthIn(nOut5_23), .SouthIn(nOut5_25), .EastIn(nOut6_24), .WestIn(nOut4_24), .ScanIn(nScanOut345), .ScanOut(nScanOut344), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_345 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_25), .NorthIn(nOut5_24), .SouthIn(nOut5_26), .EastIn(nOut6_25), .WestIn(nOut4_25), .ScanIn(nScanOut346), .ScanOut(nScanOut345), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_346 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_26), .NorthIn(nOut5_25), .SouthIn(nOut5_27), .EastIn(nOut6_26), .WestIn(nOut4_26), .ScanIn(nScanOut347), .ScanOut(nScanOut346), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_347 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_27), .NorthIn(nOut5_26), .SouthIn(nOut5_28), .EastIn(nOut6_27), .WestIn(nOut4_27), .ScanIn(nScanOut348), .ScanOut(nScanOut347), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_348 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_28), .NorthIn(nOut5_27), .SouthIn(nOut5_29), .EastIn(nOut6_28), .WestIn(nOut4_28), .ScanIn(nScanOut349), .ScanOut(nScanOut348), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_349 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_29), .NorthIn(nOut5_28), .SouthIn(nOut5_30), .EastIn(nOut6_29), .WestIn(nOut4_29), .ScanIn(nScanOut350), .ScanOut(nScanOut349), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_350 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_30), .NorthIn(nOut5_29), .SouthIn(nOut5_31), .EastIn(nOut6_30), .WestIn(nOut4_30), .ScanIn(nScanOut351), .ScanOut(nScanOut350), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_351 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_31), .NorthIn(nOut5_30), .SouthIn(nOut5_32), .EastIn(nOut6_31), .WestIn(nOut4_31), .ScanIn(nScanOut352), .ScanOut(nScanOut351), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_352 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_32), .NorthIn(nOut5_31), .SouthIn(nOut5_33), .EastIn(nOut6_32), .WestIn(nOut4_32), .ScanIn(nScanOut353), .ScanOut(nScanOut352), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_353 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_33), .NorthIn(nOut5_32), .SouthIn(nOut5_34), .EastIn(nOut6_33), .WestIn(nOut4_33), .ScanIn(nScanOut354), .ScanOut(nScanOut353), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_354 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_34), .NorthIn(nOut5_33), .SouthIn(nOut5_35), .EastIn(nOut6_34), .WestIn(nOut4_34), .ScanIn(nScanOut355), .ScanOut(nScanOut354), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_355 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_35), .NorthIn(nOut5_34), .SouthIn(nOut5_36), .EastIn(nOut6_35), .WestIn(nOut4_35), .ScanIn(nScanOut356), .ScanOut(nScanOut355), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_356 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_36), .NorthIn(nOut5_35), .SouthIn(nOut5_37), .EastIn(nOut6_36), .WestIn(nOut4_36), .ScanIn(nScanOut357), .ScanOut(nScanOut356), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_357 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_37), .NorthIn(nOut5_36), .SouthIn(nOut5_38), .EastIn(nOut6_37), .WestIn(nOut4_37), .ScanIn(nScanOut358), .ScanOut(nScanOut357), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_358 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_38), .NorthIn(nOut5_37), .SouthIn(nOut5_39), .EastIn(nOut6_38), .WestIn(nOut4_38), .ScanIn(nScanOut359), .ScanOut(nScanOut358), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_359 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_39), .NorthIn(nOut5_38), .SouthIn(nOut5_40), .EastIn(nOut6_39), .WestIn(nOut4_39), .ScanIn(nScanOut360), .ScanOut(nScanOut359), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_360 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_40), .NorthIn(nOut5_39), .SouthIn(nOut5_41), .EastIn(nOut6_40), .WestIn(nOut4_40), .ScanIn(nScanOut361), .ScanOut(nScanOut360), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_361 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_41), .NorthIn(nOut5_40), .SouthIn(nOut5_42), .EastIn(nOut6_41), .WestIn(nOut4_41), .ScanIn(nScanOut362), .ScanOut(nScanOut361), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_362 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_42), .NorthIn(nOut5_41), .SouthIn(nOut5_43), .EastIn(nOut6_42), .WestIn(nOut4_42), .ScanIn(nScanOut363), .ScanOut(nScanOut362), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_363 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_43), .NorthIn(nOut5_42), .SouthIn(nOut5_44), .EastIn(nOut6_43), .WestIn(nOut4_43), .ScanIn(nScanOut364), .ScanOut(nScanOut363), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_364 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_44), .NorthIn(nOut5_43), .SouthIn(nOut5_45), .EastIn(nOut6_44), .WestIn(nOut4_44), .ScanIn(nScanOut365), .ScanOut(nScanOut364), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_365 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_45), .NorthIn(nOut5_44), .SouthIn(nOut5_46), .EastIn(nOut6_45), .WestIn(nOut4_45), .ScanIn(nScanOut366), .ScanOut(nScanOut365), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_366 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_46), .NorthIn(nOut5_45), .SouthIn(nOut5_47), .EastIn(nOut6_46), .WestIn(nOut4_46), .ScanIn(nScanOut367), .ScanOut(nScanOut366), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_367 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_47), .NorthIn(nOut5_46), .SouthIn(nOut5_48), .EastIn(nOut6_47), .WestIn(nOut4_47), .ScanIn(nScanOut368), .ScanOut(nScanOut367), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_368 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_48), .NorthIn(nOut5_47), .SouthIn(nOut5_49), .EastIn(nOut6_48), .WestIn(nOut4_48), .ScanIn(nScanOut369), .ScanOut(nScanOut368), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_369 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_49), .NorthIn(nOut5_48), .SouthIn(nOut5_50), .EastIn(nOut6_49), .WestIn(nOut4_49), .ScanIn(nScanOut370), .ScanOut(nScanOut369), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_370 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_50), .NorthIn(nOut5_49), .SouthIn(nOut5_51), .EastIn(nOut6_50), .WestIn(nOut4_50), .ScanIn(nScanOut371), .ScanOut(nScanOut370), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_371 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_51), .NorthIn(nOut5_50), .SouthIn(nOut5_52), .EastIn(nOut6_51), .WestIn(nOut4_51), .ScanIn(nScanOut372), .ScanOut(nScanOut371), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_372 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_52), .NorthIn(nOut5_51), .SouthIn(nOut5_53), .EastIn(nOut6_52), .WestIn(nOut4_52), .ScanIn(nScanOut373), .ScanOut(nScanOut372), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_373 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_53), .NorthIn(nOut5_52), .SouthIn(nOut5_54), .EastIn(nOut6_53), .WestIn(nOut4_53), .ScanIn(nScanOut374), .ScanOut(nScanOut373), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_374 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_54), .NorthIn(nOut5_53), .SouthIn(nOut5_55), .EastIn(nOut6_54), .WestIn(nOut4_54), .ScanIn(nScanOut375), .ScanOut(nScanOut374), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_375 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_55), .NorthIn(nOut5_54), .SouthIn(nOut5_56), .EastIn(nOut6_55), .WestIn(nOut4_55), .ScanIn(nScanOut376), .ScanOut(nScanOut375), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_376 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_56), .NorthIn(nOut5_55), .SouthIn(nOut5_57), .EastIn(nOut6_56), .WestIn(nOut4_56), .ScanIn(nScanOut377), .ScanOut(nScanOut376), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_377 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_57), .NorthIn(nOut5_56), .SouthIn(nOut5_58), .EastIn(nOut6_57), .WestIn(nOut4_57), .ScanIn(nScanOut378), .ScanOut(nScanOut377), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_378 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_58), .NorthIn(nOut5_57), .SouthIn(nOut5_59), .EastIn(nOut6_58), .WestIn(nOut4_58), .ScanIn(nScanOut379), .ScanOut(nScanOut378), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_379 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_59), .NorthIn(nOut5_58), .SouthIn(nOut5_60), .EastIn(nOut6_59), .WestIn(nOut4_59), .ScanIn(nScanOut380), .ScanOut(nScanOut379), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_380 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_60), .NorthIn(nOut5_59), .SouthIn(nOut5_61), .EastIn(nOut6_60), .WestIn(nOut4_60), .ScanIn(nScanOut381), .ScanOut(nScanOut380), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_381 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_61), .NorthIn(nOut5_60), .SouthIn(nOut5_62), .EastIn(nOut6_61), .WestIn(nOut4_61), .ScanIn(nScanOut382), .ScanOut(nScanOut381), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_382 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_62), .NorthIn(nOut5_61), .SouthIn(nOut5_63), .EastIn(nOut6_62), .WestIn(nOut4_62), .ScanIn(nScanOut383), .ScanOut(nScanOut382), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_383 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_63), .ScanIn(nScanOut384), .ScanOut(nScanOut383), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_384 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_0), .ScanIn(nScanOut385), .ScanOut(nScanOut384), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_385 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_1), .NorthIn(nOut6_0), .SouthIn(nOut6_2), .EastIn(nOut7_1), .WestIn(nOut5_1), .ScanIn(nScanOut386), .ScanOut(nScanOut385), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_386 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_2), .NorthIn(nOut6_1), .SouthIn(nOut6_3), .EastIn(nOut7_2), .WestIn(nOut5_2), .ScanIn(nScanOut387), .ScanOut(nScanOut386), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_387 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_3), .NorthIn(nOut6_2), .SouthIn(nOut6_4), .EastIn(nOut7_3), .WestIn(nOut5_3), .ScanIn(nScanOut388), .ScanOut(nScanOut387), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_388 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_4), .NorthIn(nOut6_3), .SouthIn(nOut6_5), .EastIn(nOut7_4), .WestIn(nOut5_4), .ScanIn(nScanOut389), .ScanOut(nScanOut388), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_389 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_5), .NorthIn(nOut6_4), .SouthIn(nOut6_6), .EastIn(nOut7_5), .WestIn(nOut5_5), .ScanIn(nScanOut390), .ScanOut(nScanOut389), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_390 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_6), .NorthIn(nOut6_5), .SouthIn(nOut6_7), .EastIn(nOut7_6), .WestIn(nOut5_6), .ScanIn(nScanOut391), .ScanOut(nScanOut390), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_391 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_7), .NorthIn(nOut6_6), .SouthIn(nOut6_8), .EastIn(nOut7_7), .WestIn(nOut5_7), .ScanIn(nScanOut392), .ScanOut(nScanOut391), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_392 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_8), .NorthIn(nOut6_7), .SouthIn(nOut6_9), .EastIn(nOut7_8), .WestIn(nOut5_8), .ScanIn(nScanOut393), .ScanOut(nScanOut392), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_393 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_9), .NorthIn(nOut6_8), .SouthIn(nOut6_10), .EastIn(nOut7_9), .WestIn(nOut5_9), .ScanIn(nScanOut394), .ScanOut(nScanOut393), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_394 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_10), .NorthIn(nOut6_9), .SouthIn(nOut6_11), .EastIn(nOut7_10), .WestIn(nOut5_10), .ScanIn(nScanOut395), .ScanOut(nScanOut394), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_395 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_11), .NorthIn(nOut6_10), .SouthIn(nOut6_12), .EastIn(nOut7_11), .WestIn(nOut5_11), .ScanIn(nScanOut396), .ScanOut(nScanOut395), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_396 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_12), .NorthIn(nOut6_11), .SouthIn(nOut6_13), .EastIn(nOut7_12), .WestIn(nOut5_12), .ScanIn(nScanOut397), .ScanOut(nScanOut396), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_397 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_13), .NorthIn(nOut6_12), .SouthIn(nOut6_14), .EastIn(nOut7_13), .WestIn(nOut5_13), .ScanIn(nScanOut398), .ScanOut(nScanOut397), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_398 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_14), .NorthIn(nOut6_13), .SouthIn(nOut6_15), .EastIn(nOut7_14), .WestIn(nOut5_14), .ScanIn(nScanOut399), .ScanOut(nScanOut398), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_399 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_15), .NorthIn(nOut6_14), .SouthIn(nOut6_16), .EastIn(nOut7_15), .WestIn(nOut5_15), .ScanIn(nScanOut400), .ScanOut(nScanOut399), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_400 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_16), .NorthIn(nOut6_15), .SouthIn(nOut6_17), .EastIn(nOut7_16), .WestIn(nOut5_16), .ScanIn(nScanOut401), .ScanOut(nScanOut400), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_401 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_17), .NorthIn(nOut6_16), .SouthIn(nOut6_18), .EastIn(nOut7_17), .WestIn(nOut5_17), .ScanIn(nScanOut402), .ScanOut(nScanOut401), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_402 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_18), .NorthIn(nOut6_17), .SouthIn(nOut6_19), .EastIn(nOut7_18), .WestIn(nOut5_18), .ScanIn(nScanOut403), .ScanOut(nScanOut402), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_403 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_19), .NorthIn(nOut6_18), .SouthIn(nOut6_20), .EastIn(nOut7_19), .WestIn(nOut5_19), .ScanIn(nScanOut404), .ScanOut(nScanOut403), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_404 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_20), .NorthIn(nOut6_19), .SouthIn(nOut6_21), .EastIn(nOut7_20), .WestIn(nOut5_20), .ScanIn(nScanOut405), .ScanOut(nScanOut404), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_405 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_21), .NorthIn(nOut6_20), .SouthIn(nOut6_22), .EastIn(nOut7_21), .WestIn(nOut5_21), .ScanIn(nScanOut406), .ScanOut(nScanOut405), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_406 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_22), .NorthIn(nOut6_21), .SouthIn(nOut6_23), .EastIn(nOut7_22), .WestIn(nOut5_22), .ScanIn(nScanOut407), .ScanOut(nScanOut406), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_407 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_23), .NorthIn(nOut6_22), .SouthIn(nOut6_24), .EastIn(nOut7_23), .WestIn(nOut5_23), .ScanIn(nScanOut408), .ScanOut(nScanOut407), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_408 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_24), .NorthIn(nOut6_23), .SouthIn(nOut6_25), .EastIn(nOut7_24), .WestIn(nOut5_24), .ScanIn(nScanOut409), .ScanOut(nScanOut408), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_409 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_25), .NorthIn(nOut6_24), .SouthIn(nOut6_26), .EastIn(nOut7_25), .WestIn(nOut5_25), .ScanIn(nScanOut410), .ScanOut(nScanOut409), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_410 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_26), .NorthIn(nOut6_25), .SouthIn(nOut6_27), .EastIn(nOut7_26), .WestIn(nOut5_26), .ScanIn(nScanOut411), .ScanOut(nScanOut410), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_411 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_27), .NorthIn(nOut6_26), .SouthIn(nOut6_28), .EastIn(nOut7_27), .WestIn(nOut5_27), .ScanIn(nScanOut412), .ScanOut(nScanOut411), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_412 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_28), .NorthIn(nOut6_27), .SouthIn(nOut6_29), .EastIn(nOut7_28), .WestIn(nOut5_28), .ScanIn(nScanOut413), .ScanOut(nScanOut412), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_413 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_29), .NorthIn(nOut6_28), .SouthIn(nOut6_30), .EastIn(nOut7_29), .WestIn(nOut5_29), .ScanIn(nScanOut414), .ScanOut(nScanOut413), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_414 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_30), .NorthIn(nOut6_29), .SouthIn(nOut6_31), .EastIn(nOut7_30), .WestIn(nOut5_30), .ScanIn(nScanOut415), .ScanOut(nScanOut414), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_415 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_31), .NorthIn(nOut6_30), .SouthIn(nOut6_32), .EastIn(nOut7_31), .WestIn(nOut5_31), .ScanIn(nScanOut416), .ScanOut(nScanOut415), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_416 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_32), .NorthIn(nOut6_31), .SouthIn(nOut6_33), .EastIn(nOut7_32), .WestIn(nOut5_32), .ScanIn(nScanOut417), .ScanOut(nScanOut416), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_417 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_33), .NorthIn(nOut6_32), .SouthIn(nOut6_34), .EastIn(nOut7_33), .WestIn(nOut5_33), .ScanIn(nScanOut418), .ScanOut(nScanOut417), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_418 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_34), .NorthIn(nOut6_33), .SouthIn(nOut6_35), .EastIn(nOut7_34), .WestIn(nOut5_34), .ScanIn(nScanOut419), .ScanOut(nScanOut418), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_419 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_35), .NorthIn(nOut6_34), .SouthIn(nOut6_36), .EastIn(nOut7_35), .WestIn(nOut5_35), .ScanIn(nScanOut420), .ScanOut(nScanOut419), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_420 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_36), .NorthIn(nOut6_35), .SouthIn(nOut6_37), .EastIn(nOut7_36), .WestIn(nOut5_36), .ScanIn(nScanOut421), .ScanOut(nScanOut420), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_421 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_37), .NorthIn(nOut6_36), .SouthIn(nOut6_38), .EastIn(nOut7_37), .WestIn(nOut5_37), .ScanIn(nScanOut422), .ScanOut(nScanOut421), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_422 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_38), .NorthIn(nOut6_37), .SouthIn(nOut6_39), .EastIn(nOut7_38), .WestIn(nOut5_38), .ScanIn(nScanOut423), .ScanOut(nScanOut422), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_423 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_39), .NorthIn(nOut6_38), .SouthIn(nOut6_40), .EastIn(nOut7_39), .WestIn(nOut5_39), .ScanIn(nScanOut424), .ScanOut(nScanOut423), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_424 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_40), .NorthIn(nOut6_39), .SouthIn(nOut6_41), .EastIn(nOut7_40), .WestIn(nOut5_40), .ScanIn(nScanOut425), .ScanOut(nScanOut424), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_425 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_41), .NorthIn(nOut6_40), .SouthIn(nOut6_42), .EastIn(nOut7_41), .WestIn(nOut5_41), .ScanIn(nScanOut426), .ScanOut(nScanOut425), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_426 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_42), .NorthIn(nOut6_41), .SouthIn(nOut6_43), .EastIn(nOut7_42), .WestIn(nOut5_42), .ScanIn(nScanOut427), .ScanOut(nScanOut426), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_427 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_43), .NorthIn(nOut6_42), .SouthIn(nOut6_44), .EastIn(nOut7_43), .WestIn(nOut5_43), .ScanIn(nScanOut428), .ScanOut(nScanOut427), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_428 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_44), .NorthIn(nOut6_43), .SouthIn(nOut6_45), .EastIn(nOut7_44), .WestIn(nOut5_44), .ScanIn(nScanOut429), .ScanOut(nScanOut428), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_429 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_45), .NorthIn(nOut6_44), .SouthIn(nOut6_46), .EastIn(nOut7_45), .WestIn(nOut5_45), .ScanIn(nScanOut430), .ScanOut(nScanOut429), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_430 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_46), .NorthIn(nOut6_45), .SouthIn(nOut6_47), .EastIn(nOut7_46), .WestIn(nOut5_46), .ScanIn(nScanOut431), .ScanOut(nScanOut430), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_431 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_47), .NorthIn(nOut6_46), .SouthIn(nOut6_48), .EastIn(nOut7_47), .WestIn(nOut5_47), .ScanIn(nScanOut432), .ScanOut(nScanOut431), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_432 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_48), .NorthIn(nOut6_47), .SouthIn(nOut6_49), .EastIn(nOut7_48), .WestIn(nOut5_48), .ScanIn(nScanOut433), .ScanOut(nScanOut432), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_433 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_49), .NorthIn(nOut6_48), .SouthIn(nOut6_50), .EastIn(nOut7_49), .WestIn(nOut5_49), .ScanIn(nScanOut434), .ScanOut(nScanOut433), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_434 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_50), .NorthIn(nOut6_49), .SouthIn(nOut6_51), .EastIn(nOut7_50), .WestIn(nOut5_50), .ScanIn(nScanOut435), .ScanOut(nScanOut434), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_435 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_51), .NorthIn(nOut6_50), .SouthIn(nOut6_52), .EastIn(nOut7_51), .WestIn(nOut5_51), .ScanIn(nScanOut436), .ScanOut(nScanOut435), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_436 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_52), .NorthIn(nOut6_51), .SouthIn(nOut6_53), .EastIn(nOut7_52), .WestIn(nOut5_52), .ScanIn(nScanOut437), .ScanOut(nScanOut436), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_437 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_53), .NorthIn(nOut6_52), .SouthIn(nOut6_54), .EastIn(nOut7_53), .WestIn(nOut5_53), .ScanIn(nScanOut438), .ScanOut(nScanOut437), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_438 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_54), .NorthIn(nOut6_53), .SouthIn(nOut6_55), .EastIn(nOut7_54), .WestIn(nOut5_54), .ScanIn(nScanOut439), .ScanOut(nScanOut438), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_439 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_55), .NorthIn(nOut6_54), .SouthIn(nOut6_56), .EastIn(nOut7_55), .WestIn(nOut5_55), .ScanIn(nScanOut440), .ScanOut(nScanOut439), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_440 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_56), .NorthIn(nOut6_55), .SouthIn(nOut6_57), .EastIn(nOut7_56), .WestIn(nOut5_56), .ScanIn(nScanOut441), .ScanOut(nScanOut440), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_441 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_57), .NorthIn(nOut6_56), .SouthIn(nOut6_58), .EastIn(nOut7_57), .WestIn(nOut5_57), .ScanIn(nScanOut442), .ScanOut(nScanOut441), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_442 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_58), .NorthIn(nOut6_57), .SouthIn(nOut6_59), .EastIn(nOut7_58), .WestIn(nOut5_58), .ScanIn(nScanOut443), .ScanOut(nScanOut442), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_443 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_59), .NorthIn(nOut6_58), .SouthIn(nOut6_60), .EastIn(nOut7_59), .WestIn(nOut5_59), .ScanIn(nScanOut444), .ScanOut(nScanOut443), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_444 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_60), .NorthIn(nOut6_59), .SouthIn(nOut6_61), .EastIn(nOut7_60), .WestIn(nOut5_60), .ScanIn(nScanOut445), .ScanOut(nScanOut444), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_445 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_61), .NorthIn(nOut6_60), .SouthIn(nOut6_62), .EastIn(nOut7_61), .WestIn(nOut5_61), .ScanIn(nScanOut446), .ScanOut(nScanOut445), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_446 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_62), .NorthIn(nOut6_61), .SouthIn(nOut6_63), .EastIn(nOut7_62), .WestIn(nOut5_62), .ScanIn(nScanOut447), .ScanOut(nScanOut446), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_447 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_63), .ScanIn(nScanOut448), .ScanOut(nScanOut447), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_448 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_0), .ScanIn(nScanOut449), .ScanOut(nScanOut448), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_449 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_1), .NorthIn(nOut7_0), .SouthIn(nOut7_2), .EastIn(nOut8_1), .WestIn(nOut6_1), .ScanIn(nScanOut450), .ScanOut(nScanOut449), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_450 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_2), .NorthIn(nOut7_1), .SouthIn(nOut7_3), .EastIn(nOut8_2), .WestIn(nOut6_2), .ScanIn(nScanOut451), .ScanOut(nScanOut450), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_451 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_3), .NorthIn(nOut7_2), .SouthIn(nOut7_4), .EastIn(nOut8_3), .WestIn(nOut6_3), .ScanIn(nScanOut452), .ScanOut(nScanOut451), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_452 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_4), .NorthIn(nOut7_3), .SouthIn(nOut7_5), .EastIn(nOut8_4), .WestIn(nOut6_4), .ScanIn(nScanOut453), .ScanOut(nScanOut452), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_453 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_5), .NorthIn(nOut7_4), .SouthIn(nOut7_6), .EastIn(nOut8_5), .WestIn(nOut6_5), .ScanIn(nScanOut454), .ScanOut(nScanOut453), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_454 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_6), .NorthIn(nOut7_5), .SouthIn(nOut7_7), .EastIn(nOut8_6), .WestIn(nOut6_6), .ScanIn(nScanOut455), .ScanOut(nScanOut454), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_455 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_7), .NorthIn(nOut7_6), .SouthIn(nOut7_8), .EastIn(nOut8_7), .WestIn(nOut6_7), .ScanIn(nScanOut456), .ScanOut(nScanOut455), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_456 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_8), .NorthIn(nOut7_7), .SouthIn(nOut7_9), .EastIn(nOut8_8), .WestIn(nOut6_8), .ScanIn(nScanOut457), .ScanOut(nScanOut456), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_457 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_9), .NorthIn(nOut7_8), .SouthIn(nOut7_10), .EastIn(nOut8_9), .WestIn(nOut6_9), .ScanIn(nScanOut458), .ScanOut(nScanOut457), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_458 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_10), .NorthIn(nOut7_9), .SouthIn(nOut7_11), .EastIn(nOut8_10), .WestIn(nOut6_10), .ScanIn(nScanOut459), .ScanOut(nScanOut458), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_459 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_11), .NorthIn(nOut7_10), .SouthIn(nOut7_12), .EastIn(nOut8_11), .WestIn(nOut6_11), .ScanIn(nScanOut460), .ScanOut(nScanOut459), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_460 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_12), .NorthIn(nOut7_11), .SouthIn(nOut7_13), .EastIn(nOut8_12), .WestIn(nOut6_12), .ScanIn(nScanOut461), .ScanOut(nScanOut460), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_461 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_13), .NorthIn(nOut7_12), .SouthIn(nOut7_14), .EastIn(nOut8_13), .WestIn(nOut6_13), .ScanIn(nScanOut462), .ScanOut(nScanOut461), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_462 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_14), .NorthIn(nOut7_13), .SouthIn(nOut7_15), .EastIn(nOut8_14), .WestIn(nOut6_14), .ScanIn(nScanOut463), .ScanOut(nScanOut462), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_463 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_15), .NorthIn(nOut7_14), .SouthIn(nOut7_16), .EastIn(nOut8_15), .WestIn(nOut6_15), .ScanIn(nScanOut464), .ScanOut(nScanOut463), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_464 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_16), .NorthIn(nOut7_15), .SouthIn(nOut7_17), .EastIn(nOut8_16), .WestIn(nOut6_16), .ScanIn(nScanOut465), .ScanOut(nScanOut464), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_465 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_17), .NorthIn(nOut7_16), .SouthIn(nOut7_18), .EastIn(nOut8_17), .WestIn(nOut6_17), .ScanIn(nScanOut466), .ScanOut(nScanOut465), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_466 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_18), .NorthIn(nOut7_17), .SouthIn(nOut7_19), .EastIn(nOut8_18), .WestIn(nOut6_18), .ScanIn(nScanOut467), .ScanOut(nScanOut466), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_467 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_19), .NorthIn(nOut7_18), .SouthIn(nOut7_20), .EastIn(nOut8_19), .WestIn(nOut6_19), .ScanIn(nScanOut468), .ScanOut(nScanOut467), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_468 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_20), .NorthIn(nOut7_19), .SouthIn(nOut7_21), .EastIn(nOut8_20), .WestIn(nOut6_20), .ScanIn(nScanOut469), .ScanOut(nScanOut468), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_469 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_21), .NorthIn(nOut7_20), .SouthIn(nOut7_22), .EastIn(nOut8_21), .WestIn(nOut6_21), .ScanIn(nScanOut470), .ScanOut(nScanOut469), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_470 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_22), .NorthIn(nOut7_21), .SouthIn(nOut7_23), .EastIn(nOut8_22), .WestIn(nOut6_22), .ScanIn(nScanOut471), .ScanOut(nScanOut470), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_471 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_23), .NorthIn(nOut7_22), .SouthIn(nOut7_24), .EastIn(nOut8_23), .WestIn(nOut6_23), .ScanIn(nScanOut472), .ScanOut(nScanOut471), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_472 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_24), .NorthIn(nOut7_23), .SouthIn(nOut7_25), .EastIn(nOut8_24), .WestIn(nOut6_24), .ScanIn(nScanOut473), .ScanOut(nScanOut472), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_473 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_25), .NorthIn(nOut7_24), .SouthIn(nOut7_26), .EastIn(nOut8_25), .WestIn(nOut6_25), .ScanIn(nScanOut474), .ScanOut(nScanOut473), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_474 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_26), .NorthIn(nOut7_25), .SouthIn(nOut7_27), .EastIn(nOut8_26), .WestIn(nOut6_26), .ScanIn(nScanOut475), .ScanOut(nScanOut474), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_475 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_27), .NorthIn(nOut7_26), .SouthIn(nOut7_28), .EastIn(nOut8_27), .WestIn(nOut6_27), .ScanIn(nScanOut476), .ScanOut(nScanOut475), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_476 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_28), .NorthIn(nOut7_27), .SouthIn(nOut7_29), .EastIn(nOut8_28), .WestIn(nOut6_28), .ScanIn(nScanOut477), .ScanOut(nScanOut476), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_477 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_29), .NorthIn(nOut7_28), .SouthIn(nOut7_30), .EastIn(nOut8_29), .WestIn(nOut6_29), .ScanIn(nScanOut478), .ScanOut(nScanOut477), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_478 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_30), .NorthIn(nOut7_29), .SouthIn(nOut7_31), .EastIn(nOut8_30), .WestIn(nOut6_30), .ScanIn(nScanOut479), .ScanOut(nScanOut478), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_479 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_31), .NorthIn(nOut7_30), .SouthIn(nOut7_32), .EastIn(nOut8_31), .WestIn(nOut6_31), .ScanIn(nScanOut480), .ScanOut(nScanOut479), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_480 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_32), .NorthIn(nOut7_31), .SouthIn(nOut7_33), .EastIn(nOut8_32), .WestIn(nOut6_32), .ScanIn(nScanOut481), .ScanOut(nScanOut480), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_481 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_33), .NorthIn(nOut7_32), .SouthIn(nOut7_34), .EastIn(nOut8_33), .WestIn(nOut6_33), .ScanIn(nScanOut482), .ScanOut(nScanOut481), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_482 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_34), .NorthIn(nOut7_33), .SouthIn(nOut7_35), .EastIn(nOut8_34), .WestIn(nOut6_34), .ScanIn(nScanOut483), .ScanOut(nScanOut482), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_483 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_35), .NorthIn(nOut7_34), .SouthIn(nOut7_36), .EastIn(nOut8_35), .WestIn(nOut6_35), .ScanIn(nScanOut484), .ScanOut(nScanOut483), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_484 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_36), .NorthIn(nOut7_35), .SouthIn(nOut7_37), .EastIn(nOut8_36), .WestIn(nOut6_36), .ScanIn(nScanOut485), .ScanOut(nScanOut484), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_485 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_37), .NorthIn(nOut7_36), .SouthIn(nOut7_38), .EastIn(nOut8_37), .WestIn(nOut6_37), .ScanIn(nScanOut486), .ScanOut(nScanOut485), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_486 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_38), .NorthIn(nOut7_37), .SouthIn(nOut7_39), .EastIn(nOut8_38), .WestIn(nOut6_38), .ScanIn(nScanOut487), .ScanOut(nScanOut486), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_487 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_39), .NorthIn(nOut7_38), .SouthIn(nOut7_40), .EastIn(nOut8_39), .WestIn(nOut6_39), .ScanIn(nScanOut488), .ScanOut(nScanOut487), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_488 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_40), .NorthIn(nOut7_39), .SouthIn(nOut7_41), .EastIn(nOut8_40), .WestIn(nOut6_40), .ScanIn(nScanOut489), .ScanOut(nScanOut488), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_489 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_41), .NorthIn(nOut7_40), .SouthIn(nOut7_42), .EastIn(nOut8_41), .WestIn(nOut6_41), .ScanIn(nScanOut490), .ScanOut(nScanOut489), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_490 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_42), .NorthIn(nOut7_41), .SouthIn(nOut7_43), .EastIn(nOut8_42), .WestIn(nOut6_42), .ScanIn(nScanOut491), .ScanOut(nScanOut490), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_491 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_43), .NorthIn(nOut7_42), .SouthIn(nOut7_44), .EastIn(nOut8_43), .WestIn(nOut6_43), .ScanIn(nScanOut492), .ScanOut(nScanOut491), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_492 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_44), .NorthIn(nOut7_43), .SouthIn(nOut7_45), .EastIn(nOut8_44), .WestIn(nOut6_44), .ScanIn(nScanOut493), .ScanOut(nScanOut492), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_493 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_45), .NorthIn(nOut7_44), .SouthIn(nOut7_46), .EastIn(nOut8_45), .WestIn(nOut6_45), .ScanIn(nScanOut494), .ScanOut(nScanOut493), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_494 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_46), .NorthIn(nOut7_45), .SouthIn(nOut7_47), .EastIn(nOut8_46), .WestIn(nOut6_46), .ScanIn(nScanOut495), .ScanOut(nScanOut494), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_495 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_47), .NorthIn(nOut7_46), .SouthIn(nOut7_48), .EastIn(nOut8_47), .WestIn(nOut6_47), .ScanIn(nScanOut496), .ScanOut(nScanOut495), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_496 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_48), .NorthIn(nOut7_47), .SouthIn(nOut7_49), .EastIn(nOut8_48), .WestIn(nOut6_48), .ScanIn(nScanOut497), .ScanOut(nScanOut496), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_497 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_49), .NorthIn(nOut7_48), .SouthIn(nOut7_50), .EastIn(nOut8_49), .WestIn(nOut6_49), .ScanIn(nScanOut498), .ScanOut(nScanOut497), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_498 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_50), .NorthIn(nOut7_49), .SouthIn(nOut7_51), .EastIn(nOut8_50), .WestIn(nOut6_50), .ScanIn(nScanOut499), .ScanOut(nScanOut498), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_499 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_51), .NorthIn(nOut7_50), .SouthIn(nOut7_52), .EastIn(nOut8_51), .WestIn(nOut6_51), .ScanIn(nScanOut500), .ScanOut(nScanOut499), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_500 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_52), .NorthIn(nOut7_51), .SouthIn(nOut7_53), .EastIn(nOut8_52), .WestIn(nOut6_52), .ScanIn(nScanOut501), .ScanOut(nScanOut500), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_501 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_53), .NorthIn(nOut7_52), .SouthIn(nOut7_54), .EastIn(nOut8_53), .WestIn(nOut6_53), .ScanIn(nScanOut502), .ScanOut(nScanOut501), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_502 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_54), .NorthIn(nOut7_53), .SouthIn(nOut7_55), .EastIn(nOut8_54), .WestIn(nOut6_54), .ScanIn(nScanOut503), .ScanOut(nScanOut502), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_503 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_55), .NorthIn(nOut7_54), .SouthIn(nOut7_56), .EastIn(nOut8_55), .WestIn(nOut6_55), .ScanIn(nScanOut504), .ScanOut(nScanOut503), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_504 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_56), .NorthIn(nOut7_55), .SouthIn(nOut7_57), .EastIn(nOut8_56), .WestIn(nOut6_56), .ScanIn(nScanOut505), .ScanOut(nScanOut504), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_505 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_57), .NorthIn(nOut7_56), .SouthIn(nOut7_58), .EastIn(nOut8_57), .WestIn(nOut6_57), .ScanIn(nScanOut506), .ScanOut(nScanOut505), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_506 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_58), .NorthIn(nOut7_57), .SouthIn(nOut7_59), .EastIn(nOut8_58), .WestIn(nOut6_58), .ScanIn(nScanOut507), .ScanOut(nScanOut506), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_507 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_59), .NorthIn(nOut7_58), .SouthIn(nOut7_60), .EastIn(nOut8_59), .WestIn(nOut6_59), .ScanIn(nScanOut508), .ScanOut(nScanOut507), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_508 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_60), .NorthIn(nOut7_59), .SouthIn(nOut7_61), .EastIn(nOut8_60), .WestIn(nOut6_60), .ScanIn(nScanOut509), .ScanOut(nScanOut508), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_509 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_61), .NorthIn(nOut7_60), .SouthIn(nOut7_62), .EastIn(nOut8_61), .WestIn(nOut6_61), .ScanIn(nScanOut510), .ScanOut(nScanOut509), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_510 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_62), .NorthIn(nOut7_61), .SouthIn(nOut7_63), .EastIn(nOut8_62), .WestIn(nOut6_62), .ScanIn(nScanOut511), .ScanOut(nScanOut510), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_511 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_63), .ScanIn(nScanOut512), .ScanOut(nScanOut511), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_512 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut8_0), .ScanIn(nScanOut513), .ScanOut(nScanOut512), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_513 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_1), .NorthIn(nOut8_0), .SouthIn(nOut8_2), .EastIn(nOut9_1), .WestIn(nOut7_1), .ScanIn(nScanOut514), .ScanOut(nScanOut513), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_514 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_2), .NorthIn(nOut8_1), .SouthIn(nOut8_3), .EastIn(nOut9_2), .WestIn(nOut7_2), .ScanIn(nScanOut515), .ScanOut(nScanOut514), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_515 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_3), .NorthIn(nOut8_2), .SouthIn(nOut8_4), .EastIn(nOut9_3), .WestIn(nOut7_3), .ScanIn(nScanOut516), .ScanOut(nScanOut515), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_516 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_4), .NorthIn(nOut8_3), .SouthIn(nOut8_5), .EastIn(nOut9_4), .WestIn(nOut7_4), .ScanIn(nScanOut517), .ScanOut(nScanOut516), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_517 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_5), .NorthIn(nOut8_4), .SouthIn(nOut8_6), .EastIn(nOut9_5), .WestIn(nOut7_5), .ScanIn(nScanOut518), .ScanOut(nScanOut517), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_518 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_6), .NorthIn(nOut8_5), .SouthIn(nOut8_7), .EastIn(nOut9_6), .WestIn(nOut7_6), .ScanIn(nScanOut519), .ScanOut(nScanOut518), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_519 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_7), .NorthIn(nOut8_6), .SouthIn(nOut8_8), .EastIn(nOut9_7), .WestIn(nOut7_7), .ScanIn(nScanOut520), .ScanOut(nScanOut519), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_520 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_8), .NorthIn(nOut8_7), .SouthIn(nOut8_9), .EastIn(nOut9_8), .WestIn(nOut7_8), .ScanIn(nScanOut521), .ScanOut(nScanOut520), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_521 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_9), .NorthIn(nOut8_8), .SouthIn(nOut8_10), .EastIn(nOut9_9), .WestIn(nOut7_9), .ScanIn(nScanOut522), .ScanOut(nScanOut521), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_522 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_10), .NorthIn(nOut8_9), .SouthIn(nOut8_11), .EastIn(nOut9_10), .WestIn(nOut7_10), .ScanIn(nScanOut523), .ScanOut(nScanOut522), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_523 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_11), .NorthIn(nOut8_10), .SouthIn(nOut8_12), .EastIn(nOut9_11), .WestIn(nOut7_11), .ScanIn(nScanOut524), .ScanOut(nScanOut523), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_524 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_12), .NorthIn(nOut8_11), .SouthIn(nOut8_13), .EastIn(nOut9_12), .WestIn(nOut7_12), .ScanIn(nScanOut525), .ScanOut(nScanOut524), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_525 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_13), .NorthIn(nOut8_12), .SouthIn(nOut8_14), .EastIn(nOut9_13), .WestIn(nOut7_13), .ScanIn(nScanOut526), .ScanOut(nScanOut525), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_526 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_14), .NorthIn(nOut8_13), .SouthIn(nOut8_15), .EastIn(nOut9_14), .WestIn(nOut7_14), .ScanIn(nScanOut527), .ScanOut(nScanOut526), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_527 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_15), .NorthIn(nOut8_14), .SouthIn(nOut8_16), .EastIn(nOut9_15), .WestIn(nOut7_15), .ScanIn(nScanOut528), .ScanOut(nScanOut527), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_528 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_16), .NorthIn(nOut8_15), .SouthIn(nOut8_17), .EastIn(nOut9_16), .WestIn(nOut7_16), .ScanIn(nScanOut529), .ScanOut(nScanOut528), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_529 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_17), .NorthIn(nOut8_16), .SouthIn(nOut8_18), .EastIn(nOut9_17), .WestIn(nOut7_17), .ScanIn(nScanOut530), .ScanOut(nScanOut529), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_530 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_18), .NorthIn(nOut8_17), .SouthIn(nOut8_19), .EastIn(nOut9_18), .WestIn(nOut7_18), .ScanIn(nScanOut531), .ScanOut(nScanOut530), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_531 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_19), .NorthIn(nOut8_18), .SouthIn(nOut8_20), .EastIn(nOut9_19), .WestIn(nOut7_19), .ScanIn(nScanOut532), .ScanOut(nScanOut531), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_532 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_20), .NorthIn(nOut8_19), .SouthIn(nOut8_21), .EastIn(nOut9_20), .WestIn(nOut7_20), .ScanIn(nScanOut533), .ScanOut(nScanOut532), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_533 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_21), .NorthIn(nOut8_20), .SouthIn(nOut8_22), .EastIn(nOut9_21), .WestIn(nOut7_21), .ScanIn(nScanOut534), .ScanOut(nScanOut533), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_534 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_22), .NorthIn(nOut8_21), .SouthIn(nOut8_23), .EastIn(nOut9_22), .WestIn(nOut7_22), .ScanIn(nScanOut535), .ScanOut(nScanOut534), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_535 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_23), .NorthIn(nOut8_22), .SouthIn(nOut8_24), .EastIn(nOut9_23), .WestIn(nOut7_23), .ScanIn(nScanOut536), .ScanOut(nScanOut535), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_536 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_24), .NorthIn(nOut8_23), .SouthIn(nOut8_25), .EastIn(nOut9_24), .WestIn(nOut7_24), .ScanIn(nScanOut537), .ScanOut(nScanOut536), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_537 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_25), .NorthIn(nOut8_24), .SouthIn(nOut8_26), .EastIn(nOut9_25), .WestIn(nOut7_25), .ScanIn(nScanOut538), .ScanOut(nScanOut537), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_538 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_26), .NorthIn(nOut8_25), .SouthIn(nOut8_27), .EastIn(nOut9_26), .WestIn(nOut7_26), .ScanIn(nScanOut539), .ScanOut(nScanOut538), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_539 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_27), .NorthIn(nOut8_26), .SouthIn(nOut8_28), .EastIn(nOut9_27), .WestIn(nOut7_27), .ScanIn(nScanOut540), .ScanOut(nScanOut539), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_540 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_28), .NorthIn(nOut8_27), .SouthIn(nOut8_29), .EastIn(nOut9_28), .WestIn(nOut7_28), .ScanIn(nScanOut541), .ScanOut(nScanOut540), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_541 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_29), .NorthIn(nOut8_28), .SouthIn(nOut8_30), .EastIn(nOut9_29), .WestIn(nOut7_29), .ScanIn(nScanOut542), .ScanOut(nScanOut541), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_542 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_30), .NorthIn(nOut8_29), .SouthIn(nOut8_31), .EastIn(nOut9_30), .WestIn(nOut7_30), .ScanIn(nScanOut543), .ScanOut(nScanOut542), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_543 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_31), .NorthIn(nOut8_30), .SouthIn(nOut8_32), .EastIn(nOut9_31), .WestIn(nOut7_31), .ScanIn(nScanOut544), .ScanOut(nScanOut543), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_544 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_32), .NorthIn(nOut8_31), .SouthIn(nOut8_33), .EastIn(nOut9_32), .WestIn(nOut7_32), .ScanIn(nScanOut545), .ScanOut(nScanOut544), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_545 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_33), .NorthIn(nOut8_32), .SouthIn(nOut8_34), .EastIn(nOut9_33), .WestIn(nOut7_33), .ScanIn(nScanOut546), .ScanOut(nScanOut545), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_546 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_34), .NorthIn(nOut8_33), .SouthIn(nOut8_35), .EastIn(nOut9_34), .WestIn(nOut7_34), .ScanIn(nScanOut547), .ScanOut(nScanOut546), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_547 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_35), .NorthIn(nOut8_34), .SouthIn(nOut8_36), .EastIn(nOut9_35), .WestIn(nOut7_35), .ScanIn(nScanOut548), .ScanOut(nScanOut547), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_548 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_36), .NorthIn(nOut8_35), .SouthIn(nOut8_37), .EastIn(nOut9_36), .WestIn(nOut7_36), .ScanIn(nScanOut549), .ScanOut(nScanOut548), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_549 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_37), .NorthIn(nOut8_36), .SouthIn(nOut8_38), .EastIn(nOut9_37), .WestIn(nOut7_37), .ScanIn(nScanOut550), .ScanOut(nScanOut549), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_550 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_38), .NorthIn(nOut8_37), .SouthIn(nOut8_39), .EastIn(nOut9_38), .WestIn(nOut7_38), .ScanIn(nScanOut551), .ScanOut(nScanOut550), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_551 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_39), .NorthIn(nOut8_38), .SouthIn(nOut8_40), .EastIn(nOut9_39), .WestIn(nOut7_39), .ScanIn(nScanOut552), .ScanOut(nScanOut551), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_552 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_40), .NorthIn(nOut8_39), .SouthIn(nOut8_41), .EastIn(nOut9_40), .WestIn(nOut7_40), .ScanIn(nScanOut553), .ScanOut(nScanOut552), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_553 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_41), .NorthIn(nOut8_40), .SouthIn(nOut8_42), .EastIn(nOut9_41), .WestIn(nOut7_41), .ScanIn(nScanOut554), .ScanOut(nScanOut553), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_554 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_42), .NorthIn(nOut8_41), .SouthIn(nOut8_43), .EastIn(nOut9_42), .WestIn(nOut7_42), .ScanIn(nScanOut555), .ScanOut(nScanOut554), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_555 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_43), .NorthIn(nOut8_42), .SouthIn(nOut8_44), .EastIn(nOut9_43), .WestIn(nOut7_43), .ScanIn(nScanOut556), .ScanOut(nScanOut555), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_556 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_44), .NorthIn(nOut8_43), .SouthIn(nOut8_45), .EastIn(nOut9_44), .WestIn(nOut7_44), .ScanIn(nScanOut557), .ScanOut(nScanOut556), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_557 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_45), .NorthIn(nOut8_44), .SouthIn(nOut8_46), .EastIn(nOut9_45), .WestIn(nOut7_45), .ScanIn(nScanOut558), .ScanOut(nScanOut557), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_558 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_46), .NorthIn(nOut8_45), .SouthIn(nOut8_47), .EastIn(nOut9_46), .WestIn(nOut7_46), .ScanIn(nScanOut559), .ScanOut(nScanOut558), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_559 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_47), .NorthIn(nOut8_46), .SouthIn(nOut8_48), .EastIn(nOut9_47), .WestIn(nOut7_47), .ScanIn(nScanOut560), .ScanOut(nScanOut559), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_560 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_48), .NorthIn(nOut8_47), .SouthIn(nOut8_49), .EastIn(nOut9_48), .WestIn(nOut7_48), .ScanIn(nScanOut561), .ScanOut(nScanOut560), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_561 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_49), .NorthIn(nOut8_48), .SouthIn(nOut8_50), .EastIn(nOut9_49), .WestIn(nOut7_49), .ScanIn(nScanOut562), .ScanOut(nScanOut561), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_562 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_50), .NorthIn(nOut8_49), .SouthIn(nOut8_51), .EastIn(nOut9_50), .WestIn(nOut7_50), .ScanIn(nScanOut563), .ScanOut(nScanOut562), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_563 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_51), .NorthIn(nOut8_50), .SouthIn(nOut8_52), .EastIn(nOut9_51), .WestIn(nOut7_51), .ScanIn(nScanOut564), .ScanOut(nScanOut563), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_564 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_52), .NorthIn(nOut8_51), .SouthIn(nOut8_53), .EastIn(nOut9_52), .WestIn(nOut7_52), .ScanIn(nScanOut565), .ScanOut(nScanOut564), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_565 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_53), .NorthIn(nOut8_52), .SouthIn(nOut8_54), .EastIn(nOut9_53), .WestIn(nOut7_53), .ScanIn(nScanOut566), .ScanOut(nScanOut565), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_566 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_54), .NorthIn(nOut8_53), .SouthIn(nOut8_55), .EastIn(nOut9_54), .WestIn(nOut7_54), .ScanIn(nScanOut567), .ScanOut(nScanOut566), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_567 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_55), .NorthIn(nOut8_54), .SouthIn(nOut8_56), .EastIn(nOut9_55), .WestIn(nOut7_55), .ScanIn(nScanOut568), .ScanOut(nScanOut567), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_568 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_56), .NorthIn(nOut8_55), .SouthIn(nOut8_57), .EastIn(nOut9_56), .WestIn(nOut7_56), .ScanIn(nScanOut569), .ScanOut(nScanOut568), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_569 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_57), .NorthIn(nOut8_56), .SouthIn(nOut8_58), .EastIn(nOut9_57), .WestIn(nOut7_57), .ScanIn(nScanOut570), .ScanOut(nScanOut569), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_570 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_58), .NorthIn(nOut8_57), .SouthIn(nOut8_59), .EastIn(nOut9_58), .WestIn(nOut7_58), .ScanIn(nScanOut571), .ScanOut(nScanOut570), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_571 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_59), .NorthIn(nOut8_58), .SouthIn(nOut8_60), .EastIn(nOut9_59), .WestIn(nOut7_59), .ScanIn(nScanOut572), .ScanOut(nScanOut571), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_572 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_60), .NorthIn(nOut8_59), .SouthIn(nOut8_61), .EastIn(nOut9_60), .WestIn(nOut7_60), .ScanIn(nScanOut573), .ScanOut(nScanOut572), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_573 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_61), .NorthIn(nOut8_60), .SouthIn(nOut8_62), .EastIn(nOut9_61), .WestIn(nOut7_61), .ScanIn(nScanOut574), .ScanOut(nScanOut573), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_574 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_62), .NorthIn(nOut8_61), .SouthIn(nOut8_63), .EastIn(nOut9_62), .WestIn(nOut7_62), .ScanIn(nScanOut575), .ScanOut(nScanOut574), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_575 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut8_63), .ScanIn(nScanOut576), .ScanOut(nScanOut575), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_576 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut9_0), .ScanIn(nScanOut577), .ScanOut(nScanOut576), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_577 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_1), .NorthIn(nOut9_0), .SouthIn(nOut9_2), .EastIn(nOut10_1), .WestIn(nOut8_1), .ScanIn(nScanOut578), .ScanOut(nScanOut577), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_578 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_2), .NorthIn(nOut9_1), .SouthIn(nOut9_3), .EastIn(nOut10_2), .WestIn(nOut8_2), .ScanIn(nScanOut579), .ScanOut(nScanOut578), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_579 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_3), .NorthIn(nOut9_2), .SouthIn(nOut9_4), .EastIn(nOut10_3), .WestIn(nOut8_3), .ScanIn(nScanOut580), .ScanOut(nScanOut579), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_580 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_4), .NorthIn(nOut9_3), .SouthIn(nOut9_5), .EastIn(nOut10_4), .WestIn(nOut8_4), .ScanIn(nScanOut581), .ScanOut(nScanOut580), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_581 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_5), .NorthIn(nOut9_4), .SouthIn(nOut9_6), .EastIn(nOut10_5), .WestIn(nOut8_5), .ScanIn(nScanOut582), .ScanOut(nScanOut581), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_582 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_6), .NorthIn(nOut9_5), .SouthIn(nOut9_7), .EastIn(nOut10_6), .WestIn(nOut8_6), .ScanIn(nScanOut583), .ScanOut(nScanOut582), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_583 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_7), .NorthIn(nOut9_6), .SouthIn(nOut9_8), .EastIn(nOut10_7), .WestIn(nOut8_7), .ScanIn(nScanOut584), .ScanOut(nScanOut583), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_584 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_8), .NorthIn(nOut9_7), .SouthIn(nOut9_9), .EastIn(nOut10_8), .WestIn(nOut8_8), .ScanIn(nScanOut585), .ScanOut(nScanOut584), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_585 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_9), .NorthIn(nOut9_8), .SouthIn(nOut9_10), .EastIn(nOut10_9), .WestIn(nOut8_9), .ScanIn(nScanOut586), .ScanOut(nScanOut585), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_586 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_10), .NorthIn(nOut9_9), .SouthIn(nOut9_11), .EastIn(nOut10_10), .WestIn(nOut8_10), .ScanIn(nScanOut587), .ScanOut(nScanOut586), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_587 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_11), .NorthIn(nOut9_10), .SouthIn(nOut9_12), .EastIn(nOut10_11), .WestIn(nOut8_11), .ScanIn(nScanOut588), .ScanOut(nScanOut587), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_588 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_12), .NorthIn(nOut9_11), .SouthIn(nOut9_13), .EastIn(nOut10_12), .WestIn(nOut8_12), .ScanIn(nScanOut589), .ScanOut(nScanOut588), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_589 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_13), .NorthIn(nOut9_12), .SouthIn(nOut9_14), .EastIn(nOut10_13), .WestIn(nOut8_13), .ScanIn(nScanOut590), .ScanOut(nScanOut589), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_590 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_14), .NorthIn(nOut9_13), .SouthIn(nOut9_15), .EastIn(nOut10_14), .WestIn(nOut8_14), .ScanIn(nScanOut591), .ScanOut(nScanOut590), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_591 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_15), .NorthIn(nOut9_14), .SouthIn(nOut9_16), .EastIn(nOut10_15), .WestIn(nOut8_15), .ScanIn(nScanOut592), .ScanOut(nScanOut591), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_592 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_16), .NorthIn(nOut9_15), .SouthIn(nOut9_17), .EastIn(nOut10_16), .WestIn(nOut8_16), .ScanIn(nScanOut593), .ScanOut(nScanOut592), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_593 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_17), .NorthIn(nOut9_16), .SouthIn(nOut9_18), .EastIn(nOut10_17), .WestIn(nOut8_17), .ScanIn(nScanOut594), .ScanOut(nScanOut593), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_594 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_18), .NorthIn(nOut9_17), .SouthIn(nOut9_19), .EastIn(nOut10_18), .WestIn(nOut8_18), .ScanIn(nScanOut595), .ScanOut(nScanOut594), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_595 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_19), .NorthIn(nOut9_18), .SouthIn(nOut9_20), .EastIn(nOut10_19), .WestIn(nOut8_19), .ScanIn(nScanOut596), .ScanOut(nScanOut595), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_596 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_20), .NorthIn(nOut9_19), .SouthIn(nOut9_21), .EastIn(nOut10_20), .WestIn(nOut8_20), .ScanIn(nScanOut597), .ScanOut(nScanOut596), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_597 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_21), .NorthIn(nOut9_20), .SouthIn(nOut9_22), .EastIn(nOut10_21), .WestIn(nOut8_21), .ScanIn(nScanOut598), .ScanOut(nScanOut597), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_598 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_22), .NorthIn(nOut9_21), .SouthIn(nOut9_23), .EastIn(nOut10_22), .WestIn(nOut8_22), .ScanIn(nScanOut599), .ScanOut(nScanOut598), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_599 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_23), .NorthIn(nOut9_22), .SouthIn(nOut9_24), .EastIn(nOut10_23), .WestIn(nOut8_23), .ScanIn(nScanOut600), .ScanOut(nScanOut599), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_600 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_24), .NorthIn(nOut9_23), .SouthIn(nOut9_25), .EastIn(nOut10_24), .WestIn(nOut8_24), .ScanIn(nScanOut601), .ScanOut(nScanOut600), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_601 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_25), .NorthIn(nOut9_24), .SouthIn(nOut9_26), .EastIn(nOut10_25), .WestIn(nOut8_25), .ScanIn(nScanOut602), .ScanOut(nScanOut601), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_602 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_26), .NorthIn(nOut9_25), .SouthIn(nOut9_27), .EastIn(nOut10_26), .WestIn(nOut8_26), .ScanIn(nScanOut603), .ScanOut(nScanOut602), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_603 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_27), .NorthIn(nOut9_26), .SouthIn(nOut9_28), .EastIn(nOut10_27), .WestIn(nOut8_27), .ScanIn(nScanOut604), .ScanOut(nScanOut603), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_604 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_28), .NorthIn(nOut9_27), .SouthIn(nOut9_29), .EastIn(nOut10_28), .WestIn(nOut8_28), .ScanIn(nScanOut605), .ScanOut(nScanOut604), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_605 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_29), .NorthIn(nOut9_28), .SouthIn(nOut9_30), .EastIn(nOut10_29), .WestIn(nOut8_29), .ScanIn(nScanOut606), .ScanOut(nScanOut605), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_606 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_30), .NorthIn(nOut9_29), .SouthIn(nOut9_31), .EastIn(nOut10_30), .WestIn(nOut8_30), .ScanIn(nScanOut607), .ScanOut(nScanOut606), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_607 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_31), .NorthIn(nOut9_30), .SouthIn(nOut9_32), .EastIn(nOut10_31), .WestIn(nOut8_31), .ScanIn(nScanOut608), .ScanOut(nScanOut607), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_608 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_32), .NorthIn(nOut9_31), .SouthIn(nOut9_33), .EastIn(nOut10_32), .WestIn(nOut8_32), .ScanIn(nScanOut609), .ScanOut(nScanOut608), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_609 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_33), .NorthIn(nOut9_32), .SouthIn(nOut9_34), .EastIn(nOut10_33), .WestIn(nOut8_33), .ScanIn(nScanOut610), .ScanOut(nScanOut609), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_610 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_34), .NorthIn(nOut9_33), .SouthIn(nOut9_35), .EastIn(nOut10_34), .WestIn(nOut8_34), .ScanIn(nScanOut611), .ScanOut(nScanOut610), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_611 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_35), .NorthIn(nOut9_34), .SouthIn(nOut9_36), .EastIn(nOut10_35), .WestIn(nOut8_35), .ScanIn(nScanOut612), .ScanOut(nScanOut611), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_612 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_36), .NorthIn(nOut9_35), .SouthIn(nOut9_37), .EastIn(nOut10_36), .WestIn(nOut8_36), .ScanIn(nScanOut613), .ScanOut(nScanOut612), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_613 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_37), .NorthIn(nOut9_36), .SouthIn(nOut9_38), .EastIn(nOut10_37), .WestIn(nOut8_37), .ScanIn(nScanOut614), .ScanOut(nScanOut613), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_614 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_38), .NorthIn(nOut9_37), .SouthIn(nOut9_39), .EastIn(nOut10_38), .WestIn(nOut8_38), .ScanIn(nScanOut615), .ScanOut(nScanOut614), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_615 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_39), .NorthIn(nOut9_38), .SouthIn(nOut9_40), .EastIn(nOut10_39), .WestIn(nOut8_39), .ScanIn(nScanOut616), .ScanOut(nScanOut615), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_616 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_40), .NorthIn(nOut9_39), .SouthIn(nOut9_41), .EastIn(nOut10_40), .WestIn(nOut8_40), .ScanIn(nScanOut617), .ScanOut(nScanOut616), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_617 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_41), .NorthIn(nOut9_40), .SouthIn(nOut9_42), .EastIn(nOut10_41), .WestIn(nOut8_41), .ScanIn(nScanOut618), .ScanOut(nScanOut617), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_618 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_42), .NorthIn(nOut9_41), .SouthIn(nOut9_43), .EastIn(nOut10_42), .WestIn(nOut8_42), .ScanIn(nScanOut619), .ScanOut(nScanOut618), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_619 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_43), .NorthIn(nOut9_42), .SouthIn(nOut9_44), .EastIn(nOut10_43), .WestIn(nOut8_43), .ScanIn(nScanOut620), .ScanOut(nScanOut619), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_620 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_44), .NorthIn(nOut9_43), .SouthIn(nOut9_45), .EastIn(nOut10_44), .WestIn(nOut8_44), .ScanIn(nScanOut621), .ScanOut(nScanOut620), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_621 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_45), .NorthIn(nOut9_44), .SouthIn(nOut9_46), .EastIn(nOut10_45), .WestIn(nOut8_45), .ScanIn(nScanOut622), .ScanOut(nScanOut621), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_622 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_46), .NorthIn(nOut9_45), .SouthIn(nOut9_47), .EastIn(nOut10_46), .WestIn(nOut8_46), .ScanIn(nScanOut623), .ScanOut(nScanOut622), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_623 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_47), .NorthIn(nOut9_46), .SouthIn(nOut9_48), .EastIn(nOut10_47), .WestIn(nOut8_47), .ScanIn(nScanOut624), .ScanOut(nScanOut623), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_624 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_48), .NorthIn(nOut9_47), .SouthIn(nOut9_49), .EastIn(nOut10_48), .WestIn(nOut8_48), .ScanIn(nScanOut625), .ScanOut(nScanOut624), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_625 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_49), .NorthIn(nOut9_48), .SouthIn(nOut9_50), .EastIn(nOut10_49), .WestIn(nOut8_49), .ScanIn(nScanOut626), .ScanOut(nScanOut625), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_626 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_50), .NorthIn(nOut9_49), .SouthIn(nOut9_51), .EastIn(nOut10_50), .WestIn(nOut8_50), .ScanIn(nScanOut627), .ScanOut(nScanOut626), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_627 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_51), .NorthIn(nOut9_50), .SouthIn(nOut9_52), .EastIn(nOut10_51), .WestIn(nOut8_51), .ScanIn(nScanOut628), .ScanOut(nScanOut627), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_628 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_52), .NorthIn(nOut9_51), .SouthIn(nOut9_53), .EastIn(nOut10_52), .WestIn(nOut8_52), .ScanIn(nScanOut629), .ScanOut(nScanOut628), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_629 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_53), .NorthIn(nOut9_52), .SouthIn(nOut9_54), .EastIn(nOut10_53), .WestIn(nOut8_53), .ScanIn(nScanOut630), .ScanOut(nScanOut629), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_630 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_54), .NorthIn(nOut9_53), .SouthIn(nOut9_55), .EastIn(nOut10_54), .WestIn(nOut8_54), .ScanIn(nScanOut631), .ScanOut(nScanOut630), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_631 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_55), .NorthIn(nOut9_54), .SouthIn(nOut9_56), .EastIn(nOut10_55), .WestIn(nOut8_55), .ScanIn(nScanOut632), .ScanOut(nScanOut631), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_632 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_56), .NorthIn(nOut9_55), .SouthIn(nOut9_57), .EastIn(nOut10_56), .WestIn(nOut8_56), .ScanIn(nScanOut633), .ScanOut(nScanOut632), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_633 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_57), .NorthIn(nOut9_56), .SouthIn(nOut9_58), .EastIn(nOut10_57), .WestIn(nOut8_57), .ScanIn(nScanOut634), .ScanOut(nScanOut633), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_634 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_58), .NorthIn(nOut9_57), .SouthIn(nOut9_59), .EastIn(nOut10_58), .WestIn(nOut8_58), .ScanIn(nScanOut635), .ScanOut(nScanOut634), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_635 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_59), .NorthIn(nOut9_58), .SouthIn(nOut9_60), .EastIn(nOut10_59), .WestIn(nOut8_59), .ScanIn(nScanOut636), .ScanOut(nScanOut635), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_636 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_60), .NorthIn(nOut9_59), .SouthIn(nOut9_61), .EastIn(nOut10_60), .WestIn(nOut8_60), .ScanIn(nScanOut637), .ScanOut(nScanOut636), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_637 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_61), .NorthIn(nOut9_60), .SouthIn(nOut9_62), .EastIn(nOut10_61), .WestIn(nOut8_61), .ScanIn(nScanOut638), .ScanOut(nScanOut637), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_638 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_62), .NorthIn(nOut9_61), .SouthIn(nOut9_63), .EastIn(nOut10_62), .WestIn(nOut8_62), .ScanIn(nScanOut639), .ScanOut(nScanOut638), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_639 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut9_63), .ScanIn(nScanOut640), .ScanOut(nScanOut639), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_640 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut10_0), .ScanIn(nScanOut641), .ScanOut(nScanOut640), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_641 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_1), .NorthIn(nOut10_0), .SouthIn(nOut10_2), .EastIn(nOut11_1), .WestIn(nOut9_1), .ScanIn(nScanOut642), .ScanOut(nScanOut641), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_642 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_2), .NorthIn(nOut10_1), .SouthIn(nOut10_3), .EastIn(nOut11_2), .WestIn(nOut9_2), .ScanIn(nScanOut643), .ScanOut(nScanOut642), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_643 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_3), .NorthIn(nOut10_2), .SouthIn(nOut10_4), .EastIn(nOut11_3), .WestIn(nOut9_3), .ScanIn(nScanOut644), .ScanOut(nScanOut643), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_644 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_4), .NorthIn(nOut10_3), .SouthIn(nOut10_5), .EastIn(nOut11_4), .WestIn(nOut9_4), .ScanIn(nScanOut645), .ScanOut(nScanOut644), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_645 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_5), .NorthIn(nOut10_4), .SouthIn(nOut10_6), .EastIn(nOut11_5), .WestIn(nOut9_5), .ScanIn(nScanOut646), .ScanOut(nScanOut645), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_646 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_6), .NorthIn(nOut10_5), .SouthIn(nOut10_7), .EastIn(nOut11_6), .WestIn(nOut9_6), .ScanIn(nScanOut647), .ScanOut(nScanOut646), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_647 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_7), .NorthIn(nOut10_6), .SouthIn(nOut10_8), .EastIn(nOut11_7), .WestIn(nOut9_7), .ScanIn(nScanOut648), .ScanOut(nScanOut647), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_648 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_8), .NorthIn(nOut10_7), .SouthIn(nOut10_9), .EastIn(nOut11_8), .WestIn(nOut9_8), .ScanIn(nScanOut649), .ScanOut(nScanOut648), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_649 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_9), .NorthIn(nOut10_8), .SouthIn(nOut10_10), .EastIn(nOut11_9), .WestIn(nOut9_9), .ScanIn(nScanOut650), .ScanOut(nScanOut649), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_650 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_10), .NorthIn(nOut10_9), .SouthIn(nOut10_11), .EastIn(nOut11_10), .WestIn(nOut9_10), .ScanIn(nScanOut651), .ScanOut(nScanOut650), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_651 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_11), .NorthIn(nOut10_10), .SouthIn(nOut10_12), .EastIn(nOut11_11), .WestIn(nOut9_11), .ScanIn(nScanOut652), .ScanOut(nScanOut651), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_652 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_12), .NorthIn(nOut10_11), .SouthIn(nOut10_13), .EastIn(nOut11_12), .WestIn(nOut9_12), .ScanIn(nScanOut653), .ScanOut(nScanOut652), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_653 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_13), .NorthIn(nOut10_12), .SouthIn(nOut10_14), .EastIn(nOut11_13), .WestIn(nOut9_13), .ScanIn(nScanOut654), .ScanOut(nScanOut653), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_654 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_14), .NorthIn(nOut10_13), .SouthIn(nOut10_15), .EastIn(nOut11_14), .WestIn(nOut9_14), .ScanIn(nScanOut655), .ScanOut(nScanOut654), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_655 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_15), .NorthIn(nOut10_14), .SouthIn(nOut10_16), .EastIn(nOut11_15), .WestIn(nOut9_15), .ScanIn(nScanOut656), .ScanOut(nScanOut655), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_656 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_16), .NorthIn(nOut10_15), .SouthIn(nOut10_17), .EastIn(nOut11_16), .WestIn(nOut9_16), .ScanIn(nScanOut657), .ScanOut(nScanOut656), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_657 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_17), .NorthIn(nOut10_16), .SouthIn(nOut10_18), .EastIn(nOut11_17), .WestIn(nOut9_17), .ScanIn(nScanOut658), .ScanOut(nScanOut657), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_658 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_18), .NorthIn(nOut10_17), .SouthIn(nOut10_19), .EastIn(nOut11_18), .WestIn(nOut9_18), .ScanIn(nScanOut659), .ScanOut(nScanOut658), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_659 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_19), .NorthIn(nOut10_18), .SouthIn(nOut10_20), .EastIn(nOut11_19), .WestIn(nOut9_19), .ScanIn(nScanOut660), .ScanOut(nScanOut659), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_660 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_20), .NorthIn(nOut10_19), .SouthIn(nOut10_21), .EastIn(nOut11_20), .WestIn(nOut9_20), .ScanIn(nScanOut661), .ScanOut(nScanOut660), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_661 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_21), .NorthIn(nOut10_20), .SouthIn(nOut10_22), .EastIn(nOut11_21), .WestIn(nOut9_21), .ScanIn(nScanOut662), .ScanOut(nScanOut661), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_662 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_22), .NorthIn(nOut10_21), .SouthIn(nOut10_23), .EastIn(nOut11_22), .WestIn(nOut9_22), .ScanIn(nScanOut663), .ScanOut(nScanOut662), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_663 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_23), .NorthIn(nOut10_22), .SouthIn(nOut10_24), .EastIn(nOut11_23), .WestIn(nOut9_23), .ScanIn(nScanOut664), .ScanOut(nScanOut663), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_664 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_24), .NorthIn(nOut10_23), .SouthIn(nOut10_25), .EastIn(nOut11_24), .WestIn(nOut9_24), .ScanIn(nScanOut665), .ScanOut(nScanOut664), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_665 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_25), .NorthIn(nOut10_24), .SouthIn(nOut10_26), .EastIn(nOut11_25), .WestIn(nOut9_25), .ScanIn(nScanOut666), .ScanOut(nScanOut665), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_666 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_26), .NorthIn(nOut10_25), .SouthIn(nOut10_27), .EastIn(nOut11_26), .WestIn(nOut9_26), .ScanIn(nScanOut667), .ScanOut(nScanOut666), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_667 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_27), .NorthIn(nOut10_26), .SouthIn(nOut10_28), .EastIn(nOut11_27), .WestIn(nOut9_27), .ScanIn(nScanOut668), .ScanOut(nScanOut667), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_668 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_28), .NorthIn(nOut10_27), .SouthIn(nOut10_29), .EastIn(nOut11_28), .WestIn(nOut9_28), .ScanIn(nScanOut669), .ScanOut(nScanOut668), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_669 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_29), .NorthIn(nOut10_28), .SouthIn(nOut10_30), .EastIn(nOut11_29), .WestIn(nOut9_29), .ScanIn(nScanOut670), .ScanOut(nScanOut669), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_670 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_30), .NorthIn(nOut10_29), .SouthIn(nOut10_31), .EastIn(nOut11_30), .WestIn(nOut9_30), .ScanIn(nScanOut671), .ScanOut(nScanOut670), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_671 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_31), .NorthIn(nOut10_30), .SouthIn(nOut10_32), .EastIn(nOut11_31), .WestIn(nOut9_31), .ScanIn(nScanOut672), .ScanOut(nScanOut671), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_672 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_32), .NorthIn(nOut10_31), .SouthIn(nOut10_33), .EastIn(nOut11_32), .WestIn(nOut9_32), .ScanIn(nScanOut673), .ScanOut(nScanOut672), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_673 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_33), .NorthIn(nOut10_32), .SouthIn(nOut10_34), .EastIn(nOut11_33), .WestIn(nOut9_33), .ScanIn(nScanOut674), .ScanOut(nScanOut673), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_674 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_34), .NorthIn(nOut10_33), .SouthIn(nOut10_35), .EastIn(nOut11_34), .WestIn(nOut9_34), .ScanIn(nScanOut675), .ScanOut(nScanOut674), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_675 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_35), .NorthIn(nOut10_34), .SouthIn(nOut10_36), .EastIn(nOut11_35), .WestIn(nOut9_35), .ScanIn(nScanOut676), .ScanOut(nScanOut675), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_676 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_36), .NorthIn(nOut10_35), .SouthIn(nOut10_37), .EastIn(nOut11_36), .WestIn(nOut9_36), .ScanIn(nScanOut677), .ScanOut(nScanOut676), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_677 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_37), .NorthIn(nOut10_36), .SouthIn(nOut10_38), .EastIn(nOut11_37), .WestIn(nOut9_37), .ScanIn(nScanOut678), .ScanOut(nScanOut677), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_678 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_38), .NorthIn(nOut10_37), .SouthIn(nOut10_39), .EastIn(nOut11_38), .WestIn(nOut9_38), .ScanIn(nScanOut679), .ScanOut(nScanOut678), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_679 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_39), .NorthIn(nOut10_38), .SouthIn(nOut10_40), .EastIn(nOut11_39), .WestIn(nOut9_39), .ScanIn(nScanOut680), .ScanOut(nScanOut679), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_680 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_40), .NorthIn(nOut10_39), .SouthIn(nOut10_41), .EastIn(nOut11_40), .WestIn(nOut9_40), .ScanIn(nScanOut681), .ScanOut(nScanOut680), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_681 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_41), .NorthIn(nOut10_40), .SouthIn(nOut10_42), .EastIn(nOut11_41), .WestIn(nOut9_41), .ScanIn(nScanOut682), .ScanOut(nScanOut681), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_682 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_42), .NorthIn(nOut10_41), .SouthIn(nOut10_43), .EastIn(nOut11_42), .WestIn(nOut9_42), .ScanIn(nScanOut683), .ScanOut(nScanOut682), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_683 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_43), .NorthIn(nOut10_42), .SouthIn(nOut10_44), .EastIn(nOut11_43), .WestIn(nOut9_43), .ScanIn(nScanOut684), .ScanOut(nScanOut683), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_684 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_44), .NorthIn(nOut10_43), .SouthIn(nOut10_45), .EastIn(nOut11_44), .WestIn(nOut9_44), .ScanIn(nScanOut685), .ScanOut(nScanOut684), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_685 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_45), .NorthIn(nOut10_44), .SouthIn(nOut10_46), .EastIn(nOut11_45), .WestIn(nOut9_45), .ScanIn(nScanOut686), .ScanOut(nScanOut685), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_686 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_46), .NorthIn(nOut10_45), .SouthIn(nOut10_47), .EastIn(nOut11_46), .WestIn(nOut9_46), .ScanIn(nScanOut687), .ScanOut(nScanOut686), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_687 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_47), .NorthIn(nOut10_46), .SouthIn(nOut10_48), .EastIn(nOut11_47), .WestIn(nOut9_47), .ScanIn(nScanOut688), .ScanOut(nScanOut687), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_688 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_48), .NorthIn(nOut10_47), .SouthIn(nOut10_49), .EastIn(nOut11_48), .WestIn(nOut9_48), .ScanIn(nScanOut689), .ScanOut(nScanOut688), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_689 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_49), .NorthIn(nOut10_48), .SouthIn(nOut10_50), .EastIn(nOut11_49), .WestIn(nOut9_49), .ScanIn(nScanOut690), .ScanOut(nScanOut689), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_690 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_50), .NorthIn(nOut10_49), .SouthIn(nOut10_51), .EastIn(nOut11_50), .WestIn(nOut9_50), .ScanIn(nScanOut691), .ScanOut(nScanOut690), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_691 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_51), .NorthIn(nOut10_50), .SouthIn(nOut10_52), .EastIn(nOut11_51), .WestIn(nOut9_51), .ScanIn(nScanOut692), .ScanOut(nScanOut691), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_692 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_52), .NorthIn(nOut10_51), .SouthIn(nOut10_53), .EastIn(nOut11_52), .WestIn(nOut9_52), .ScanIn(nScanOut693), .ScanOut(nScanOut692), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_693 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_53), .NorthIn(nOut10_52), .SouthIn(nOut10_54), .EastIn(nOut11_53), .WestIn(nOut9_53), .ScanIn(nScanOut694), .ScanOut(nScanOut693), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_694 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_54), .NorthIn(nOut10_53), .SouthIn(nOut10_55), .EastIn(nOut11_54), .WestIn(nOut9_54), .ScanIn(nScanOut695), .ScanOut(nScanOut694), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_695 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_55), .NorthIn(nOut10_54), .SouthIn(nOut10_56), .EastIn(nOut11_55), .WestIn(nOut9_55), .ScanIn(nScanOut696), .ScanOut(nScanOut695), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_696 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_56), .NorthIn(nOut10_55), .SouthIn(nOut10_57), .EastIn(nOut11_56), .WestIn(nOut9_56), .ScanIn(nScanOut697), .ScanOut(nScanOut696), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_697 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_57), .NorthIn(nOut10_56), .SouthIn(nOut10_58), .EastIn(nOut11_57), .WestIn(nOut9_57), .ScanIn(nScanOut698), .ScanOut(nScanOut697), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_698 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_58), .NorthIn(nOut10_57), .SouthIn(nOut10_59), .EastIn(nOut11_58), .WestIn(nOut9_58), .ScanIn(nScanOut699), .ScanOut(nScanOut698), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_699 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_59), .NorthIn(nOut10_58), .SouthIn(nOut10_60), .EastIn(nOut11_59), .WestIn(nOut9_59), .ScanIn(nScanOut700), .ScanOut(nScanOut699), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_700 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_60), .NorthIn(nOut10_59), .SouthIn(nOut10_61), .EastIn(nOut11_60), .WestIn(nOut9_60), .ScanIn(nScanOut701), .ScanOut(nScanOut700), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_701 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_61), .NorthIn(nOut10_60), .SouthIn(nOut10_62), .EastIn(nOut11_61), .WestIn(nOut9_61), .ScanIn(nScanOut702), .ScanOut(nScanOut701), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_702 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_62), .NorthIn(nOut10_61), .SouthIn(nOut10_63), .EastIn(nOut11_62), .WestIn(nOut9_62), .ScanIn(nScanOut703), .ScanOut(nScanOut702), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_703 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut10_63), .ScanIn(nScanOut704), .ScanOut(nScanOut703), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_704 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut11_0), .ScanIn(nScanOut705), .ScanOut(nScanOut704), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_705 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_1), .NorthIn(nOut11_0), .SouthIn(nOut11_2), .EastIn(nOut12_1), .WestIn(nOut10_1), .ScanIn(nScanOut706), .ScanOut(nScanOut705), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_706 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_2), .NorthIn(nOut11_1), .SouthIn(nOut11_3), .EastIn(nOut12_2), .WestIn(nOut10_2), .ScanIn(nScanOut707), .ScanOut(nScanOut706), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_707 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_3), .NorthIn(nOut11_2), .SouthIn(nOut11_4), .EastIn(nOut12_3), .WestIn(nOut10_3), .ScanIn(nScanOut708), .ScanOut(nScanOut707), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_708 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_4), .NorthIn(nOut11_3), .SouthIn(nOut11_5), .EastIn(nOut12_4), .WestIn(nOut10_4), .ScanIn(nScanOut709), .ScanOut(nScanOut708), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_709 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_5), .NorthIn(nOut11_4), .SouthIn(nOut11_6), .EastIn(nOut12_5), .WestIn(nOut10_5), .ScanIn(nScanOut710), .ScanOut(nScanOut709), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_710 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_6), .NorthIn(nOut11_5), .SouthIn(nOut11_7), .EastIn(nOut12_6), .WestIn(nOut10_6), .ScanIn(nScanOut711), .ScanOut(nScanOut710), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_711 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_7), .NorthIn(nOut11_6), .SouthIn(nOut11_8), .EastIn(nOut12_7), .WestIn(nOut10_7), .ScanIn(nScanOut712), .ScanOut(nScanOut711), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_712 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_8), .NorthIn(nOut11_7), .SouthIn(nOut11_9), .EastIn(nOut12_8), .WestIn(nOut10_8), .ScanIn(nScanOut713), .ScanOut(nScanOut712), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_713 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_9), .NorthIn(nOut11_8), .SouthIn(nOut11_10), .EastIn(nOut12_9), .WestIn(nOut10_9), .ScanIn(nScanOut714), .ScanOut(nScanOut713), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_714 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_10), .NorthIn(nOut11_9), .SouthIn(nOut11_11), .EastIn(nOut12_10), .WestIn(nOut10_10), .ScanIn(nScanOut715), .ScanOut(nScanOut714), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_715 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_11), .NorthIn(nOut11_10), .SouthIn(nOut11_12), .EastIn(nOut12_11), .WestIn(nOut10_11), .ScanIn(nScanOut716), .ScanOut(nScanOut715), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_716 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_12), .NorthIn(nOut11_11), .SouthIn(nOut11_13), .EastIn(nOut12_12), .WestIn(nOut10_12), .ScanIn(nScanOut717), .ScanOut(nScanOut716), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_717 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_13), .NorthIn(nOut11_12), .SouthIn(nOut11_14), .EastIn(nOut12_13), .WestIn(nOut10_13), .ScanIn(nScanOut718), .ScanOut(nScanOut717), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_718 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_14), .NorthIn(nOut11_13), .SouthIn(nOut11_15), .EastIn(nOut12_14), .WestIn(nOut10_14), .ScanIn(nScanOut719), .ScanOut(nScanOut718), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_719 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_15), .NorthIn(nOut11_14), .SouthIn(nOut11_16), .EastIn(nOut12_15), .WestIn(nOut10_15), .ScanIn(nScanOut720), .ScanOut(nScanOut719), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_720 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_16), .NorthIn(nOut11_15), .SouthIn(nOut11_17), .EastIn(nOut12_16), .WestIn(nOut10_16), .ScanIn(nScanOut721), .ScanOut(nScanOut720), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_721 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_17), .NorthIn(nOut11_16), .SouthIn(nOut11_18), .EastIn(nOut12_17), .WestIn(nOut10_17), .ScanIn(nScanOut722), .ScanOut(nScanOut721), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_722 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_18), .NorthIn(nOut11_17), .SouthIn(nOut11_19), .EastIn(nOut12_18), .WestIn(nOut10_18), .ScanIn(nScanOut723), .ScanOut(nScanOut722), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_723 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_19), .NorthIn(nOut11_18), .SouthIn(nOut11_20), .EastIn(nOut12_19), .WestIn(nOut10_19), .ScanIn(nScanOut724), .ScanOut(nScanOut723), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_724 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_20), .NorthIn(nOut11_19), .SouthIn(nOut11_21), .EastIn(nOut12_20), .WestIn(nOut10_20), .ScanIn(nScanOut725), .ScanOut(nScanOut724), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_725 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_21), .NorthIn(nOut11_20), .SouthIn(nOut11_22), .EastIn(nOut12_21), .WestIn(nOut10_21), .ScanIn(nScanOut726), .ScanOut(nScanOut725), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_726 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_22), .NorthIn(nOut11_21), .SouthIn(nOut11_23), .EastIn(nOut12_22), .WestIn(nOut10_22), .ScanIn(nScanOut727), .ScanOut(nScanOut726), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_727 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_23), .NorthIn(nOut11_22), .SouthIn(nOut11_24), .EastIn(nOut12_23), .WestIn(nOut10_23), .ScanIn(nScanOut728), .ScanOut(nScanOut727), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_728 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_24), .NorthIn(nOut11_23), .SouthIn(nOut11_25), .EastIn(nOut12_24), .WestIn(nOut10_24), .ScanIn(nScanOut729), .ScanOut(nScanOut728), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_729 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_25), .NorthIn(nOut11_24), .SouthIn(nOut11_26), .EastIn(nOut12_25), .WestIn(nOut10_25), .ScanIn(nScanOut730), .ScanOut(nScanOut729), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_730 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_26), .NorthIn(nOut11_25), .SouthIn(nOut11_27), .EastIn(nOut12_26), .WestIn(nOut10_26), .ScanIn(nScanOut731), .ScanOut(nScanOut730), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_731 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_27), .NorthIn(nOut11_26), .SouthIn(nOut11_28), .EastIn(nOut12_27), .WestIn(nOut10_27), .ScanIn(nScanOut732), .ScanOut(nScanOut731), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_732 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_28), .NorthIn(nOut11_27), .SouthIn(nOut11_29), .EastIn(nOut12_28), .WestIn(nOut10_28), .ScanIn(nScanOut733), .ScanOut(nScanOut732), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_733 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_29), .NorthIn(nOut11_28), .SouthIn(nOut11_30), .EastIn(nOut12_29), .WestIn(nOut10_29), .ScanIn(nScanOut734), .ScanOut(nScanOut733), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_734 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_30), .NorthIn(nOut11_29), .SouthIn(nOut11_31), .EastIn(nOut12_30), .WestIn(nOut10_30), .ScanIn(nScanOut735), .ScanOut(nScanOut734), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_735 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_31), .NorthIn(nOut11_30), .SouthIn(nOut11_32), .EastIn(nOut12_31), .WestIn(nOut10_31), .ScanIn(nScanOut736), .ScanOut(nScanOut735), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_736 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_32), .NorthIn(nOut11_31), .SouthIn(nOut11_33), .EastIn(nOut12_32), .WestIn(nOut10_32), .ScanIn(nScanOut737), .ScanOut(nScanOut736), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_737 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_33), .NorthIn(nOut11_32), .SouthIn(nOut11_34), .EastIn(nOut12_33), .WestIn(nOut10_33), .ScanIn(nScanOut738), .ScanOut(nScanOut737), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_738 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_34), .NorthIn(nOut11_33), .SouthIn(nOut11_35), .EastIn(nOut12_34), .WestIn(nOut10_34), .ScanIn(nScanOut739), .ScanOut(nScanOut738), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_739 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_35), .NorthIn(nOut11_34), .SouthIn(nOut11_36), .EastIn(nOut12_35), .WestIn(nOut10_35), .ScanIn(nScanOut740), .ScanOut(nScanOut739), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_740 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_36), .NorthIn(nOut11_35), .SouthIn(nOut11_37), .EastIn(nOut12_36), .WestIn(nOut10_36), .ScanIn(nScanOut741), .ScanOut(nScanOut740), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_741 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_37), .NorthIn(nOut11_36), .SouthIn(nOut11_38), .EastIn(nOut12_37), .WestIn(nOut10_37), .ScanIn(nScanOut742), .ScanOut(nScanOut741), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_742 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_38), .NorthIn(nOut11_37), .SouthIn(nOut11_39), .EastIn(nOut12_38), .WestIn(nOut10_38), .ScanIn(nScanOut743), .ScanOut(nScanOut742), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_743 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_39), .NorthIn(nOut11_38), .SouthIn(nOut11_40), .EastIn(nOut12_39), .WestIn(nOut10_39), .ScanIn(nScanOut744), .ScanOut(nScanOut743), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_744 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_40), .NorthIn(nOut11_39), .SouthIn(nOut11_41), .EastIn(nOut12_40), .WestIn(nOut10_40), .ScanIn(nScanOut745), .ScanOut(nScanOut744), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_745 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_41), .NorthIn(nOut11_40), .SouthIn(nOut11_42), .EastIn(nOut12_41), .WestIn(nOut10_41), .ScanIn(nScanOut746), .ScanOut(nScanOut745), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_746 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_42), .NorthIn(nOut11_41), .SouthIn(nOut11_43), .EastIn(nOut12_42), .WestIn(nOut10_42), .ScanIn(nScanOut747), .ScanOut(nScanOut746), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_747 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_43), .NorthIn(nOut11_42), .SouthIn(nOut11_44), .EastIn(nOut12_43), .WestIn(nOut10_43), .ScanIn(nScanOut748), .ScanOut(nScanOut747), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_748 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_44), .NorthIn(nOut11_43), .SouthIn(nOut11_45), .EastIn(nOut12_44), .WestIn(nOut10_44), .ScanIn(nScanOut749), .ScanOut(nScanOut748), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_749 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_45), .NorthIn(nOut11_44), .SouthIn(nOut11_46), .EastIn(nOut12_45), .WestIn(nOut10_45), .ScanIn(nScanOut750), .ScanOut(nScanOut749), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_750 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_46), .NorthIn(nOut11_45), .SouthIn(nOut11_47), .EastIn(nOut12_46), .WestIn(nOut10_46), .ScanIn(nScanOut751), .ScanOut(nScanOut750), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_751 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_47), .NorthIn(nOut11_46), .SouthIn(nOut11_48), .EastIn(nOut12_47), .WestIn(nOut10_47), .ScanIn(nScanOut752), .ScanOut(nScanOut751), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_752 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_48), .NorthIn(nOut11_47), .SouthIn(nOut11_49), .EastIn(nOut12_48), .WestIn(nOut10_48), .ScanIn(nScanOut753), .ScanOut(nScanOut752), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_753 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_49), .NorthIn(nOut11_48), .SouthIn(nOut11_50), .EastIn(nOut12_49), .WestIn(nOut10_49), .ScanIn(nScanOut754), .ScanOut(nScanOut753), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_754 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_50), .NorthIn(nOut11_49), .SouthIn(nOut11_51), .EastIn(nOut12_50), .WestIn(nOut10_50), .ScanIn(nScanOut755), .ScanOut(nScanOut754), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_755 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_51), .NorthIn(nOut11_50), .SouthIn(nOut11_52), .EastIn(nOut12_51), .WestIn(nOut10_51), .ScanIn(nScanOut756), .ScanOut(nScanOut755), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_756 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_52), .NorthIn(nOut11_51), .SouthIn(nOut11_53), .EastIn(nOut12_52), .WestIn(nOut10_52), .ScanIn(nScanOut757), .ScanOut(nScanOut756), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_757 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_53), .NorthIn(nOut11_52), .SouthIn(nOut11_54), .EastIn(nOut12_53), .WestIn(nOut10_53), .ScanIn(nScanOut758), .ScanOut(nScanOut757), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_758 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_54), .NorthIn(nOut11_53), .SouthIn(nOut11_55), .EastIn(nOut12_54), .WestIn(nOut10_54), .ScanIn(nScanOut759), .ScanOut(nScanOut758), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_759 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_55), .NorthIn(nOut11_54), .SouthIn(nOut11_56), .EastIn(nOut12_55), .WestIn(nOut10_55), .ScanIn(nScanOut760), .ScanOut(nScanOut759), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_760 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_56), .NorthIn(nOut11_55), .SouthIn(nOut11_57), .EastIn(nOut12_56), .WestIn(nOut10_56), .ScanIn(nScanOut761), .ScanOut(nScanOut760), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_761 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_57), .NorthIn(nOut11_56), .SouthIn(nOut11_58), .EastIn(nOut12_57), .WestIn(nOut10_57), .ScanIn(nScanOut762), .ScanOut(nScanOut761), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_762 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_58), .NorthIn(nOut11_57), .SouthIn(nOut11_59), .EastIn(nOut12_58), .WestIn(nOut10_58), .ScanIn(nScanOut763), .ScanOut(nScanOut762), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_763 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_59), .NorthIn(nOut11_58), .SouthIn(nOut11_60), .EastIn(nOut12_59), .WestIn(nOut10_59), .ScanIn(nScanOut764), .ScanOut(nScanOut763), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_764 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_60), .NorthIn(nOut11_59), .SouthIn(nOut11_61), .EastIn(nOut12_60), .WestIn(nOut10_60), .ScanIn(nScanOut765), .ScanOut(nScanOut764), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_765 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_61), .NorthIn(nOut11_60), .SouthIn(nOut11_62), .EastIn(nOut12_61), .WestIn(nOut10_61), .ScanIn(nScanOut766), .ScanOut(nScanOut765), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_766 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_62), .NorthIn(nOut11_61), .SouthIn(nOut11_63), .EastIn(nOut12_62), .WestIn(nOut10_62), .ScanIn(nScanOut767), .ScanOut(nScanOut766), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_767 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut11_63), .ScanIn(nScanOut768), .ScanOut(nScanOut767), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_768 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut12_0), .ScanIn(nScanOut769), .ScanOut(nScanOut768), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_769 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_1), .NorthIn(nOut12_0), .SouthIn(nOut12_2), .EastIn(nOut13_1), .WestIn(nOut11_1), .ScanIn(nScanOut770), .ScanOut(nScanOut769), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_770 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_2), .NorthIn(nOut12_1), .SouthIn(nOut12_3), .EastIn(nOut13_2), .WestIn(nOut11_2), .ScanIn(nScanOut771), .ScanOut(nScanOut770), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_771 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_3), .NorthIn(nOut12_2), .SouthIn(nOut12_4), .EastIn(nOut13_3), .WestIn(nOut11_3), .ScanIn(nScanOut772), .ScanOut(nScanOut771), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_772 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_4), .NorthIn(nOut12_3), .SouthIn(nOut12_5), .EastIn(nOut13_4), .WestIn(nOut11_4), .ScanIn(nScanOut773), .ScanOut(nScanOut772), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_773 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_5), .NorthIn(nOut12_4), .SouthIn(nOut12_6), .EastIn(nOut13_5), .WestIn(nOut11_5), .ScanIn(nScanOut774), .ScanOut(nScanOut773), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_774 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_6), .NorthIn(nOut12_5), .SouthIn(nOut12_7), .EastIn(nOut13_6), .WestIn(nOut11_6), .ScanIn(nScanOut775), .ScanOut(nScanOut774), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_775 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_7), .NorthIn(nOut12_6), .SouthIn(nOut12_8), .EastIn(nOut13_7), .WestIn(nOut11_7), .ScanIn(nScanOut776), .ScanOut(nScanOut775), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_776 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_8), .NorthIn(nOut12_7), .SouthIn(nOut12_9), .EastIn(nOut13_8), .WestIn(nOut11_8), .ScanIn(nScanOut777), .ScanOut(nScanOut776), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_777 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_9), .NorthIn(nOut12_8), .SouthIn(nOut12_10), .EastIn(nOut13_9), .WestIn(nOut11_9), .ScanIn(nScanOut778), .ScanOut(nScanOut777), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_778 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_10), .NorthIn(nOut12_9), .SouthIn(nOut12_11), .EastIn(nOut13_10), .WestIn(nOut11_10), .ScanIn(nScanOut779), .ScanOut(nScanOut778), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_779 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_11), .NorthIn(nOut12_10), .SouthIn(nOut12_12), .EastIn(nOut13_11), .WestIn(nOut11_11), .ScanIn(nScanOut780), .ScanOut(nScanOut779), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_780 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_12), .NorthIn(nOut12_11), .SouthIn(nOut12_13), .EastIn(nOut13_12), .WestIn(nOut11_12), .ScanIn(nScanOut781), .ScanOut(nScanOut780), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_781 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_13), .NorthIn(nOut12_12), .SouthIn(nOut12_14), .EastIn(nOut13_13), .WestIn(nOut11_13), .ScanIn(nScanOut782), .ScanOut(nScanOut781), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_782 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_14), .NorthIn(nOut12_13), .SouthIn(nOut12_15), .EastIn(nOut13_14), .WestIn(nOut11_14), .ScanIn(nScanOut783), .ScanOut(nScanOut782), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_783 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_15), .NorthIn(nOut12_14), .SouthIn(nOut12_16), .EastIn(nOut13_15), .WestIn(nOut11_15), .ScanIn(nScanOut784), .ScanOut(nScanOut783), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_784 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_16), .NorthIn(nOut12_15), .SouthIn(nOut12_17), .EastIn(nOut13_16), .WestIn(nOut11_16), .ScanIn(nScanOut785), .ScanOut(nScanOut784), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_785 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_17), .NorthIn(nOut12_16), .SouthIn(nOut12_18), .EastIn(nOut13_17), .WestIn(nOut11_17), .ScanIn(nScanOut786), .ScanOut(nScanOut785), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_786 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_18), .NorthIn(nOut12_17), .SouthIn(nOut12_19), .EastIn(nOut13_18), .WestIn(nOut11_18), .ScanIn(nScanOut787), .ScanOut(nScanOut786), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_787 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_19), .NorthIn(nOut12_18), .SouthIn(nOut12_20), .EastIn(nOut13_19), .WestIn(nOut11_19), .ScanIn(nScanOut788), .ScanOut(nScanOut787), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_788 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_20), .NorthIn(nOut12_19), .SouthIn(nOut12_21), .EastIn(nOut13_20), .WestIn(nOut11_20), .ScanIn(nScanOut789), .ScanOut(nScanOut788), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_789 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_21), .NorthIn(nOut12_20), .SouthIn(nOut12_22), .EastIn(nOut13_21), .WestIn(nOut11_21), .ScanIn(nScanOut790), .ScanOut(nScanOut789), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_790 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_22), .NorthIn(nOut12_21), .SouthIn(nOut12_23), .EastIn(nOut13_22), .WestIn(nOut11_22), .ScanIn(nScanOut791), .ScanOut(nScanOut790), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_791 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_23), .NorthIn(nOut12_22), .SouthIn(nOut12_24), .EastIn(nOut13_23), .WestIn(nOut11_23), .ScanIn(nScanOut792), .ScanOut(nScanOut791), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_792 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_24), .NorthIn(nOut12_23), .SouthIn(nOut12_25), .EastIn(nOut13_24), .WestIn(nOut11_24), .ScanIn(nScanOut793), .ScanOut(nScanOut792), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_793 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_25), .NorthIn(nOut12_24), .SouthIn(nOut12_26), .EastIn(nOut13_25), .WestIn(nOut11_25), .ScanIn(nScanOut794), .ScanOut(nScanOut793), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_794 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_26), .NorthIn(nOut12_25), .SouthIn(nOut12_27), .EastIn(nOut13_26), .WestIn(nOut11_26), .ScanIn(nScanOut795), .ScanOut(nScanOut794), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_795 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_27), .NorthIn(nOut12_26), .SouthIn(nOut12_28), .EastIn(nOut13_27), .WestIn(nOut11_27), .ScanIn(nScanOut796), .ScanOut(nScanOut795), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_796 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_28), .NorthIn(nOut12_27), .SouthIn(nOut12_29), .EastIn(nOut13_28), .WestIn(nOut11_28), .ScanIn(nScanOut797), .ScanOut(nScanOut796), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_797 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_29), .NorthIn(nOut12_28), .SouthIn(nOut12_30), .EastIn(nOut13_29), .WestIn(nOut11_29), .ScanIn(nScanOut798), .ScanOut(nScanOut797), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_798 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_30), .NorthIn(nOut12_29), .SouthIn(nOut12_31), .EastIn(nOut13_30), .WestIn(nOut11_30), .ScanIn(nScanOut799), .ScanOut(nScanOut798), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_799 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_31), .NorthIn(nOut12_30), .SouthIn(nOut12_32), .EastIn(nOut13_31), .WestIn(nOut11_31), .ScanIn(nScanOut800), .ScanOut(nScanOut799), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_800 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_32), .NorthIn(nOut12_31), .SouthIn(nOut12_33), .EastIn(nOut13_32), .WestIn(nOut11_32), .ScanIn(nScanOut801), .ScanOut(nScanOut800), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_801 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_33), .NorthIn(nOut12_32), .SouthIn(nOut12_34), .EastIn(nOut13_33), .WestIn(nOut11_33), .ScanIn(nScanOut802), .ScanOut(nScanOut801), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_802 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_34), .NorthIn(nOut12_33), .SouthIn(nOut12_35), .EastIn(nOut13_34), .WestIn(nOut11_34), .ScanIn(nScanOut803), .ScanOut(nScanOut802), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_803 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_35), .NorthIn(nOut12_34), .SouthIn(nOut12_36), .EastIn(nOut13_35), .WestIn(nOut11_35), .ScanIn(nScanOut804), .ScanOut(nScanOut803), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_804 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_36), .NorthIn(nOut12_35), .SouthIn(nOut12_37), .EastIn(nOut13_36), .WestIn(nOut11_36), .ScanIn(nScanOut805), .ScanOut(nScanOut804), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_805 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_37), .NorthIn(nOut12_36), .SouthIn(nOut12_38), .EastIn(nOut13_37), .WestIn(nOut11_37), .ScanIn(nScanOut806), .ScanOut(nScanOut805), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_806 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_38), .NorthIn(nOut12_37), .SouthIn(nOut12_39), .EastIn(nOut13_38), .WestIn(nOut11_38), .ScanIn(nScanOut807), .ScanOut(nScanOut806), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_807 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_39), .NorthIn(nOut12_38), .SouthIn(nOut12_40), .EastIn(nOut13_39), .WestIn(nOut11_39), .ScanIn(nScanOut808), .ScanOut(nScanOut807), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_808 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_40), .NorthIn(nOut12_39), .SouthIn(nOut12_41), .EastIn(nOut13_40), .WestIn(nOut11_40), .ScanIn(nScanOut809), .ScanOut(nScanOut808), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_809 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_41), .NorthIn(nOut12_40), .SouthIn(nOut12_42), .EastIn(nOut13_41), .WestIn(nOut11_41), .ScanIn(nScanOut810), .ScanOut(nScanOut809), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_810 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_42), .NorthIn(nOut12_41), .SouthIn(nOut12_43), .EastIn(nOut13_42), .WestIn(nOut11_42), .ScanIn(nScanOut811), .ScanOut(nScanOut810), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_811 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_43), .NorthIn(nOut12_42), .SouthIn(nOut12_44), .EastIn(nOut13_43), .WestIn(nOut11_43), .ScanIn(nScanOut812), .ScanOut(nScanOut811), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_812 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_44), .NorthIn(nOut12_43), .SouthIn(nOut12_45), .EastIn(nOut13_44), .WestIn(nOut11_44), .ScanIn(nScanOut813), .ScanOut(nScanOut812), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_813 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_45), .NorthIn(nOut12_44), .SouthIn(nOut12_46), .EastIn(nOut13_45), .WestIn(nOut11_45), .ScanIn(nScanOut814), .ScanOut(nScanOut813), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_814 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_46), .NorthIn(nOut12_45), .SouthIn(nOut12_47), .EastIn(nOut13_46), .WestIn(nOut11_46), .ScanIn(nScanOut815), .ScanOut(nScanOut814), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_815 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_47), .NorthIn(nOut12_46), .SouthIn(nOut12_48), .EastIn(nOut13_47), .WestIn(nOut11_47), .ScanIn(nScanOut816), .ScanOut(nScanOut815), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_816 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_48), .NorthIn(nOut12_47), .SouthIn(nOut12_49), .EastIn(nOut13_48), .WestIn(nOut11_48), .ScanIn(nScanOut817), .ScanOut(nScanOut816), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_817 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_49), .NorthIn(nOut12_48), .SouthIn(nOut12_50), .EastIn(nOut13_49), .WestIn(nOut11_49), .ScanIn(nScanOut818), .ScanOut(nScanOut817), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_818 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_50), .NorthIn(nOut12_49), .SouthIn(nOut12_51), .EastIn(nOut13_50), .WestIn(nOut11_50), .ScanIn(nScanOut819), .ScanOut(nScanOut818), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_819 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_51), .NorthIn(nOut12_50), .SouthIn(nOut12_52), .EastIn(nOut13_51), .WestIn(nOut11_51), .ScanIn(nScanOut820), .ScanOut(nScanOut819), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_820 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_52), .NorthIn(nOut12_51), .SouthIn(nOut12_53), .EastIn(nOut13_52), .WestIn(nOut11_52), .ScanIn(nScanOut821), .ScanOut(nScanOut820), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_821 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_53), .NorthIn(nOut12_52), .SouthIn(nOut12_54), .EastIn(nOut13_53), .WestIn(nOut11_53), .ScanIn(nScanOut822), .ScanOut(nScanOut821), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_822 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_54), .NorthIn(nOut12_53), .SouthIn(nOut12_55), .EastIn(nOut13_54), .WestIn(nOut11_54), .ScanIn(nScanOut823), .ScanOut(nScanOut822), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_823 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_55), .NorthIn(nOut12_54), .SouthIn(nOut12_56), .EastIn(nOut13_55), .WestIn(nOut11_55), .ScanIn(nScanOut824), .ScanOut(nScanOut823), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_824 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_56), .NorthIn(nOut12_55), .SouthIn(nOut12_57), .EastIn(nOut13_56), .WestIn(nOut11_56), .ScanIn(nScanOut825), .ScanOut(nScanOut824), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_825 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_57), .NorthIn(nOut12_56), .SouthIn(nOut12_58), .EastIn(nOut13_57), .WestIn(nOut11_57), .ScanIn(nScanOut826), .ScanOut(nScanOut825), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_826 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_58), .NorthIn(nOut12_57), .SouthIn(nOut12_59), .EastIn(nOut13_58), .WestIn(nOut11_58), .ScanIn(nScanOut827), .ScanOut(nScanOut826), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_827 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_59), .NorthIn(nOut12_58), .SouthIn(nOut12_60), .EastIn(nOut13_59), .WestIn(nOut11_59), .ScanIn(nScanOut828), .ScanOut(nScanOut827), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_828 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_60), .NorthIn(nOut12_59), .SouthIn(nOut12_61), .EastIn(nOut13_60), .WestIn(nOut11_60), .ScanIn(nScanOut829), .ScanOut(nScanOut828), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_829 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_61), .NorthIn(nOut12_60), .SouthIn(nOut12_62), .EastIn(nOut13_61), .WestIn(nOut11_61), .ScanIn(nScanOut830), .ScanOut(nScanOut829), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_830 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_62), .NorthIn(nOut12_61), .SouthIn(nOut12_63), .EastIn(nOut13_62), .WestIn(nOut11_62), .ScanIn(nScanOut831), .ScanOut(nScanOut830), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_831 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut12_63), .ScanIn(nScanOut832), .ScanOut(nScanOut831), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_832 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut13_0), .ScanIn(nScanOut833), .ScanOut(nScanOut832), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_833 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_1), .NorthIn(nOut13_0), .SouthIn(nOut13_2), .EastIn(nOut14_1), .WestIn(nOut12_1), .ScanIn(nScanOut834), .ScanOut(nScanOut833), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_834 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_2), .NorthIn(nOut13_1), .SouthIn(nOut13_3), .EastIn(nOut14_2), .WestIn(nOut12_2), .ScanIn(nScanOut835), .ScanOut(nScanOut834), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_835 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_3), .NorthIn(nOut13_2), .SouthIn(nOut13_4), .EastIn(nOut14_3), .WestIn(nOut12_3), .ScanIn(nScanOut836), .ScanOut(nScanOut835), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_836 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_4), .NorthIn(nOut13_3), .SouthIn(nOut13_5), .EastIn(nOut14_4), .WestIn(nOut12_4), .ScanIn(nScanOut837), .ScanOut(nScanOut836), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_837 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_5), .NorthIn(nOut13_4), .SouthIn(nOut13_6), .EastIn(nOut14_5), .WestIn(nOut12_5), .ScanIn(nScanOut838), .ScanOut(nScanOut837), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_838 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_6), .NorthIn(nOut13_5), .SouthIn(nOut13_7), .EastIn(nOut14_6), .WestIn(nOut12_6), .ScanIn(nScanOut839), .ScanOut(nScanOut838), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_839 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_7), .NorthIn(nOut13_6), .SouthIn(nOut13_8), .EastIn(nOut14_7), .WestIn(nOut12_7), .ScanIn(nScanOut840), .ScanOut(nScanOut839), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_840 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_8), .NorthIn(nOut13_7), .SouthIn(nOut13_9), .EastIn(nOut14_8), .WestIn(nOut12_8), .ScanIn(nScanOut841), .ScanOut(nScanOut840), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_841 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_9), .NorthIn(nOut13_8), .SouthIn(nOut13_10), .EastIn(nOut14_9), .WestIn(nOut12_9), .ScanIn(nScanOut842), .ScanOut(nScanOut841), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_842 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_10), .NorthIn(nOut13_9), .SouthIn(nOut13_11), .EastIn(nOut14_10), .WestIn(nOut12_10), .ScanIn(nScanOut843), .ScanOut(nScanOut842), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_843 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_11), .NorthIn(nOut13_10), .SouthIn(nOut13_12), .EastIn(nOut14_11), .WestIn(nOut12_11), .ScanIn(nScanOut844), .ScanOut(nScanOut843), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_844 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_12), .NorthIn(nOut13_11), .SouthIn(nOut13_13), .EastIn(nOut14_12), .WestIn(nOut12_12), .ScanIn(nScanOut845), .ScanOut(nScanOut844), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_845 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_13), .NorthIn(nOut13_12), .SouthIn(nOut13_14), .EastIn(nOut14_13), .WestIn(nOut12_13), .ScanIn(nScanOut846), .ScanOut(nScanOut845), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_846 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_14), .NorthIn(nOut13_13), .SouthIn(nOut13_15), .EastIn(nOut14_14), .WestIn(nOut12_14), .ScanIn(nScanOut847), .ScanOut(nScanOut846), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_847 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_15), .NorthIn(nOut13_14), .SouthIn(nOut13_16), .EastIn(nOut14_15), .WestIn(nOut12_15), .ScanIn(nScanOut848), .ScanOut(nScanOut847), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_848 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_16), .NorthIn(nOut13_15), .SouthIn(nOut13_17), .EastIn(nOut14_16), .WestIn(nOut12_16), .ScanIn(nScanOut849), .ScanOut(nScanOut848), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_849 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_17), .NorthIn(nOut13_16), .SouthIn(nOut13_18), .EastIn(nOut14_17), .WestIn(nOut12_17), .ScanIn(nScanOut850), .ScanOut(nScanOut849), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_850 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_18), .NorthIn(nOut13_17), .SouthIn(nOut13_19), .EastIn(nOut14_18), .WestIn(nOut12_18), .ScanIn(nScanOut851), .ScanOut(nScanOut850), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_851 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_19), .NorthIn(nOut13_18), .SouthIn(nOut13_20), .EastIn(nOut14_19), .WestIn(nOut12_19), .ScanIn(nScanOut852), .ScanOut(nScanOut851), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_852 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_20), .NorthIn(nOut13_19), .SouthIn(nOut13_21), .EastIn(nOut14_20), .WestIn(nOut12_20), .ScanIn(nScanOut853), .ScanOut(nScanOut852), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_853 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_21), .NorthIn(nOut13_20), .SouthIn(nOut13_22), .EastIn(nOut14_21), .WestIn(nOut12_21), .ScanIn(nScanOut854), .ScanOut(nScanOut853), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_854 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_22), .NorthIn(nOut13_21), .SouthIn(nOut13_23), .EastIn(nOut14_22), .WestIn(nOut12_22), .ScanIn(nScanOut855), .ScanOut(nScanOut854), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_855 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_23), .NorthIn(nOut13_22), .SouthIn(nOut13_24), .EastIn(nOut14_23), .WestIn(nOut12_23), .ScanIn(nScanOut856), .ScanOut(nScanOut855), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_856 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_24), .NorthIn(nOut13_23), .SouthIn(nOut13_25), .EastIn(nOut14_24), .WestIn(nOut12_24), .ScanIn(nScanOut857), .ScanOut(nScanOut856), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_857 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_25), .NorthIn(nOut13_24), .SouthIn(nOut13_26), .EastIn(nOut14_25), .WestIn(nOut12_25), .ScanIn(nScanOut858), .ScanOut(nScanOut857), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_858 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_26), .NorthIn(nOut13_25), .SouthIn(nOut13_27), .EastIn(nOut14_26), .WestIn(nOut12_26), .ScanIn(nScanOut859), .ScanOut(nScanOut858), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_859 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_27), .NorthIn(nOut13_26), .SouthIn(nOut13_28), .EastIn(nOut14_27), .WestIn(nOut12_27), .ScanIn(nScanOut860), .ScanOut(nScanOut859), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_860 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_28), .NorthIn(nOut13_27), .SouthIn(nOut13_29), .EastIn(nOut14_28), .WestIn(nOut12_28), .ScanIn(nScanOut861), .ScanOut(nScanOut860), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_861 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_29), .NorthIn(nOut13_28), .SouthIn(nOut13_30), .EastIn(nOut14_29), .WestIn(nOut12_29), .ScanIn(nScanOut862), .ScanOut(nScanOut861), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_862 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_30), .NorthIn(nOut13_29), .SouthIn(nOut13_31), .EastIn(nOut14_30), .WestIn(nOut12_30), .ScanIn(nScanOut863), .ScanOut(nScanOut862), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_863 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_31), .NorthIn(nOut13_30), .SouthIn(nOut13_32), .EastIn(nOut14_31), .WestIn(nOut12_31), .ScanIn(nScanOut864), .ScanOut(nScanOut863), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_864 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_32), .NorthIn(nOut13_31), .SouthIn(nOut13_33), .EastIn(nOut14_32), .WestIn(nOut12_32), .ScanIn(nScanOut865), .ScanOut(nScanOut864), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_865 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_33), .NorthIn(nOut13_32), .SouthIn(nOut13_34), .EastIn(nOut14_33), .WestIn(nOut12_33), .ScanIn(nScanOut866), .ScanOut(nScanOut865), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_866 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_34), .NorthIn(nOut13_33), .SouthIn(nOut13_35), .EastIn(nOut14_34), .WestIn(nOut12_34), .ScanIn(nScanOut867), .ScanOut(nScanOut866), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_867 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_35), .NorthIn(nOut13_34), .SouthIn(nOut13_36), .EastIn(nOut14_35), .WestIn(nOut12_35), .ScanIn(nScanOut868), .ScanOut(nScanOut867), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_868 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_36), .NorthIn(nOut13_35), .SouthIn(nOut13_37), .EastIn(nOut14_36), .WestIn(nOut12_36), .ScanIn(nScanOut869), .ScanOut(nScanOut868), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_869 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_37), .NorthIn(nOut13_36), .SouthIn(nOut13_38), .EastIn(nOut14_37), .WestIn(nOut12_37), .ScanIn(nScanOut870), .ScanOut(nScanOut869), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_870 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_38), .NorthIn(nOut13_37), .SouthIn(nOut13_39), .EastIn(nOut14_38), .WestIn(nOut12_38), .ScanIn(nScanOut871), .ScanOut(nScanOut870), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_871 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_39), .NorthIn(nOut13_38), .SouthIn(nOut13_40), .EastIn(nOut14_39), .WestIn(nOut12_39), .ScanIn(nScanOut872), .ScanOut(nScanOut871), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_872 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_40), .NorthIn(nOut13_39), .SouthIn(nOut13_41), .EastIn(nOut14_40), .WestIn(nOut12_40), .ScanIn(nScanOut873), .ScanOut(nScanOut872), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_873 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_41), .NorthIn(nOut13_40), .SouthIn(nOut13_42), .EastIn(nOut14_41), .WestIn(nOut12_41), .ScanIn(nScanOut874), .ScanOut(nScanOut873), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_874 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_42), .NorthIn(nOut13_41), .SouthIn(nOut13_43), .EastIn(nOut14_42), .WestIn(nOut12_42), .ScanIn(nScanOut875), .ScanOut(nScanOut874), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_875 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_43), .NorthIn(nOut13_42), .SouthIn(nOut13_44), .EastIn(nOut14_43), .WestIn(nOut12_43), .ScanIn(nScanOut876), .ScanOut(nScanOut875), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_876 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_44), .NorthIn(nOut13_43), .SouthIn(nOut13_45), .EastIn(nOut14_44), .WestIn(nOut12_44), .ScanIn(nScanOut877), .ScanOut(nScanOut876), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_877 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_45), .NorthIn(nOut13_44), .SouthIn(nOut13_46), .EastIn(nOut14_45), .WestIn(nOut12_45), .ScanIn(nScanOut878), .ScanOut(nScanOut877), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_878 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_46), .NorthIn(nOut13_45), .SouthIn(nOut13_47), .EastIn(nOut14_46), .WestIn(nOut12_46), .ScanIn(nScanOut879), .ScanOut(nScanOut878), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_879 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_47), .NorthIn(nOut13_46), .SouthIn(nOut13_48), .EastIn(nOut14_47), .WestIn(nOut12_47), .ScanIn(nScanOut880), .ScanOut(nScanOut879), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_880 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_48), .NorthIn(nOut13_47), .SouthIn(nOut13_49), .EastIn(nOut14_48), .WestIn(nOut12_48), .ScanIn(nScanOut881), .ScanOut(nScanOut880), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_881 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_49), .NorthIn(nOut13_48), .SouthIn(nOut13_50), .EastIn(nOut14_49), .WestIn(nOut12_49), .ScanIn(nScanOut882), .ScanOut(nScanOut881), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_882 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_50), .NorthIn(nOut13_49), .SouthIn(nOut13_51), .EastIn(nOut14_50), .WestIn(nOut12_50), .ScanIn(nScanOut883), .ScanOut(nScanOut882), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_883 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_51), .NorthIn(nOut13_50), .SouthIn(nOut13_52), .EastIn(nOut14_51), .WestIn(nOut12_51), .ScanIn(nScanOut884), .ScanOut(nScanOut883), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_884 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_52), .NorthIn(nOut13_51), .SouthIn(nOut13_53), .EastIn(nOut14_52), .WestIn(nOut12_52), .ScanIn(nScanOut885), .ScanOut(nScanOut884), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_885 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_53), .NorthIn(nOut13_52), .SouthIn(nOut13_54), .EastIn(nOut14_53), .WestIn(nOut12_53), .ScanIn(nScanOut886), .ScanOut(nScanOut885), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_886 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_54), .NorthIn(nOut13_53), .SouthIn(nOut13_55), .EastIn(nOut14_54), .WestIn(nOut12_54), .ScanIn(nScanOut887), .ScanOut(nScanOut886), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_887 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_55), .NorthIn(nOut13_54), .SouthIn(nOut13_56), .EastIn(nOut14_55), .WestIn(nOut12_55), .ScanIn(nScanOut888), .ScanOut(nScanOut887), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_888 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_56), .NorthIn(nOut13_55), .SouthIn(nOut13_57), .EastIn(nOut14_56), .WestIn(nOut12_56), .ScanIn(nScanOut889), .ScanOut(nScanOut888), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_889 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_57), .NorthIn(nOut13_56), .SouthIn(nOut13_58), .EastIn(nOut14_57), .WestIn(nOut12_57), .ScanIn(nScanOut890), .ScanOut(nScanOut889), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_890 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_58), .NorthIn(nOut13_57), .SouthIn(nOut13_59), .EastIn(nOut14_58), .WestIn(nOut12_58), .ScanIn(nScanOut891), .ScanOut(nScanOut890), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_891 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_59), .NorthIn(nOut13_58), .SouthIn(nOut13_60), .EastIn(nOut14_59), .WestIn(nOut12_59), .ScanIn(nScanOut892), .ScanOut(nScanOut891), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_892 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_60), .NorthIn(nOut13_59), .SouthIn(nOut13_61), .EastIn(nOut14_60), .WestIn(nOut12_60), .ScanIn(nScanOut893), .ScanOut(nScanOut892), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_893 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_61), .NorthIn(nOut13_60), .SouthIn(nOut13_62), .EastIn(nOut14_61), .WestIn(nOut12_61), .ScanIn(nScanOut894), .ScanOut(nScanOut893), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_894 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_62), .NorthIn(nOut13_61), .SouthIn(nOut13_63), .EastIn(nOut14_62), .WestIn(nOut12_62), .ScanIn(nScanOut895), .ScanOut(nScanOut894), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_895 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut13_63), .ScanIn(nScanOut896), .ScanOut(nScanOut895), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_896 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut14_0), .ScanIn(nScanOut897), .ScanOut(nScanOut896), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_897 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_1), .NorthIn(nOut14_0), .SouthIn(nOut14_2), .EastIn(nOut15_1), .WestIn(nOut13_1), .ScanIn(nScanOut898), .ScanOut(nScanOut897), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_898 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_2), .NorthIn(nOut14_1), .SouthIn(nOut14_3), .EastIn(nOut15_2), .WestIn(nOut13_2), .ScanIn(nScanOut899), .ScanOut(nScanOut898), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_899 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_3), .NorthIn(nOut14_2), .SouthIn(nOut14_4), .EastIn(nOut15_3), .WestIn(nOut13_3), .ScanIn(nScanOut900), .ScanOut(nScanOut899), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_900 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_4), .NorthIn(nOut14_3), .SouthIn(nOut14_5), .EastIn(nOut15_4), .WestIn(nOut13_4), .ScanIn(nScanOut901), .ScanOut(nScanOut900), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_901 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_5), .NorthIn(nOut14_4), .SouthIn(nOut14_6), .EastIn(nOut15_5), .WestIn(nOut13_5), .ScanIn(nScanOut902), .ScanOut(nScanOut901), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_902 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_6), .NorthIn(nOut14_5), .SouthIn(nOut14_7), .EastIn(nOut15_6), .WestIn(nOut13_6), .ScanIn(nScanOut903), .ScanOut(nScanOut902), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_903 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_7), .NorthIn(nOut14_6), .SouthIn(nOut14_8), .EastIn(nOut15_7), .WestIn(nOut13_7), .ScanIn(nScanOut904), .ScanOut(nScanOut903), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_904 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_8), .NorthIn(nOut14_7), .SouthIn(nOut14_9), .EastIn(nOut15_8), .WestIn(nOut13_8), .ScanIn(nScanOut905), .ScanOut(nScanOut904), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_905 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_9), .NorthIn(nOut14_8), .SouthIn(nOut14_10), .EastIn(nOut15_9), .WestIn(nOut13_9), .ScanIn(nScanOut906), .ScanOut(nScanOut905), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_906 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_10), .NorthIn(nOut14_9), .SouthIn(nOut14_11), .EastIn(nOut15_10), .WestIn(nOut13_10), .ScanIn(nScanOut907), .ScanOut(nScanOut906), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_907 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_11), .NorthIn(nOut14_10), .SouthIn(nOut14_12), .EastIn(nOut15_11), .WestIn(nOut13_11), .ScanIn(nScanOut908), .ScanOut(nScanOut907), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_908 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_12), .NorthIn(nOut14_11), .SouthIn(nOut14_13), .EastIn(nOut15_12), .WestIn(nOut13_12), .ScanIn(nScanOut909), .ScanOut(nScanOut908), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_909 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_13), .NorthIn(nOut14_12), .SouthIn(nOut14_14), .EastIn(nOut15_13), .WestIn(nOut13_13), .ScanIn(nScanOut910), .ScanOut(nScanOut909), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_910 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_14), .NorthIn(nOut14_13), .SouthIn(nOut14_15), .EastIn(nOut15_14), .WestIn(nOut13_14), .ScanIn(nScanOut911), .ScanOut(nScanOut910), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_911 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_15), .NorthIn(nOut14_14), .SouthIn(nOut14_16), .EastIn(nOut15_15), .WestIn(nOut13_15), .ScanIn(nScanOut912), .ScanOut(nScanOut911), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_912 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_16), .NorthIn(nOut14_15), .SouthIn(nOut14_17), .EastIn(nOut15_16), .WestIn(nOut13_16), .ScanIn(nScanOut913), .ScanOut(nScanOut912), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_913 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_17), .NorthIn(nOut14_16), .SouthIn(nOut14_18), .EastIn(nOut15_17), .WestIn(nOut13_17), .ScanIn(nScanOut914), .ScanOut(nScanOut913), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_914 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_18), .NorthIn(nOut14_17), .SouthIn(nOut14_19), .EastIn(nOut15_18), .WestIn(nOut13_18), .ScanIn(nScanOut915), .ScanOut(nScanOut914), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_915 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_19), .NorthIn(nOut14_18), .SouthIn(nOut14_20), .EastIn(nOut15_19), .WestIn(nOut13_19), .ScanIn(nScanOut916), .ScanOut(nScanOut915), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_916 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_20), .NorthIn(nOut14_19), .SouthIn(nOut14_21), .EastIn(nOut15_20), .WestIn(nOut13_20), .ScanIn(nScanOut917), .ScanOut(nScanOut916), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_917 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_21), .NorthIn(nOut14_20), .SouthIn(nOut14_22), .EastIn(nOut15_21), .WestIn(nOut13_21), .ScanIn(nScanOut918), .ScanOut(nScanOut917), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_918 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_22), .NorthIn(nOut14_21), .SouthIn(nOut14_23), .EastIn(nOut15_22), .WestIn(nOut13_22), .ScanIn(nScanOut919), .ScanOut(nScanOut918), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_919 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_23), .NorthIn(nOut14_22), .SouthIn(nOut14_24), .EastIn(nOut15_23), .WestIn(nOut13_23), .ScanIn(nScanOut920), .ScanOut(nScanOut919), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_920 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_24), .NorthIn(nOut14_23), .SouthIn(nOut14_25), .EastIn(nOut15_24), .WestIn(nOut13_24), .ScanIn(nScanOut921), .ScanOut(nScanOut920), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_921 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_25), .NorthIn(nOut14_24), .SouthIn(nOut14_26), .EastIn(nOut15_25), .WestIn(nOut13_25), .ScanIn(nScanOut922), .ScanOut(nScanOut921), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_922 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_26), .NorthIn(nOut14_25), .SouthIn(nOut14_27), .EastIn(nOut15_26), .WestIn(nOut13_26), .ScanIn(nScanOut923), .ScanOut(nScanOut922), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_923 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_27), .NorthIn(nOut14_26), .SouthIn(nOut14_28), .EastIn(nOut15_27), .WestIn(nOut13_27), .ScanIn(nScanOut924), .ScanOut(nScanOut923), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_924 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_28), .NorthIn(nOut14_27), .SouthIn(nOut14_29), .EastIn(nOut15_28), .WestIn(nOut13_28), .ScanIn(nScanOut925), .ScanOut(nScanOut924), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_925 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_29), .NorthIn(nOut14_28), .SouthIn(nOut14_30), .EastIn(nOut15_29), .WestIn(nOut13_29), .ScanIn(nScanOut926), .ScanOut(nScanOut925), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_926 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_30), .NorthIn(nOut14_29), .SouthIn(nOut14_31), .EastIn(nOut15_30), .WestIn(nOut13_30), .ScanIn(nScanOut927), .ScanOut(nScanOut926), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_927 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_31), .NorthIn(nOut14_30), .SouthIn(nOut14_32), .EastIn(nOut15_31), .WestIn(nOut13_31), .ScanIn(nScanOut928), .ScanOut(nScanOut927), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_928 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_32), .NorthIn(nOut14_31), .SouthIn(nOut14_33), .EastIn(nOut15_32), .WestIn(nOut13_32), .ScanIn(nScanOut929), .ScanOut(nScanOut928), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_929 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_33), .NorthIn(nOut14_32), .SouthIn(nOut14_34), .EastIn(nOut15_33), .WestIn(nOut13_33), .ScanIn(nScanOut930), .ScanOut(nScanOut929), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_930 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_34), .NorthIn(nOut14_33), .SouthIn(nOut14_35), .EastIn(nOut15_34), .WestIn(nOut13_34), .ScanIn(nScanOut931), .ScanOut(nScanOut930), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_931 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_35), .NorthIn(nOut14_34), .SouthIn(nOut14_36), .EastIn(nOut15_35), .WestIn(nOut13_35), .ScanIn(nScanOut932), .ScanOut(nScanOut931), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_932 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_36), .NorthIn(nOut14_35), .SouthIn(nOut14_37), .EastIn(nOut15_36), .WestIn(nOut13_36), .ScanIn(nScanOut933), .ScanOut(nScanOut932), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_933 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_37), .NorthIn(nOut14_36), .SouthIn(nOut14_38), .EastIn(nOut15_37), .WestIn(nOut13_37), .ScanIn(nScanOut934), .ScanOut(nScanOut933), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_934 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_38), .NorthIn(nOut14_37), .SouthIn(nOut14_39), .EastIn(nOut15_38), .WestIn(nOut13_38), .ScanIn(nScanOut935), .ScanOut(nScanOut934), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_935 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_39), .NorthIn(nOut14_38), .SouthIn(nOut14_40), .EastIn(nOut15_39), .WestIn(nOut13_39), .ScanIn(nScanOut936), .ScanOut(nScanOut935), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_936 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_40), .NorthIn(nOut14_39), .SouthIn(nOut14_41), .EastIn(nOut15_40), .WestIn(nOut13_40), .ScanIn(nScanOut937), .ScanOut(nScanOut936), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_937 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_41), .NorthIn(nOut14_40), .SouthIn(nOut14_42), .EastIn(nOut15_41), .WestIn(nOut13_41), .ScanIn(nScanOut938), .ScanOut(nScanOut937), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_938 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_42), .NorthIn(nOut14_41), .SouthIn(nOut14_43), .EastIn(nOut15_42), .WestIn(nOut13_42), .ScanIn(nScanOut939), .ScanOut(nScanOut938), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_939 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_43), .NorthIn(nOut14_42), .SouthIn(nOut14_44), .EastIn(nOut15_43), .WestIn(nOut13_43), .ScanIn(nScanOut940), .ScanOut(nScanOut939), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_940 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_44), .NorthIn(nOut14_43), .SouthIn(nOut14_45), .EastIn(nOut15_44), .WestIn(nOut13_44), .ScanIn(nScanOut941), .ScanOut(nScanOut940), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_941 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_45), .NorthIn(nOut14_44), .SouthIn(nOut14_46), .EastIn(nOut15_45), .WestIn(nOut13_45), .ScanIn(nScanOut942), .ScanOut(nScanOut941), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_942 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_46), .NorthIn(nOut14_45), .SouthIn(nOut14_47), .EastIn(nOut15_46), .WestIn(nOut13_46), .ScanIn(nScanOut943), .ScanOut(nScanOut942), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_943 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_47), .NorthIn(nOut14_46), .SouthIn(nOut14_48), .EastIn(nOut15_47), .WestIn(nOut13_47), .ScanIn(nScanOut944), .ScanOut(nScanOut943), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_944 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_48), .NorthIn(nOut14_47), .SouthIn(nOut14_49), .EastIn(nOut15_48), .WestIn(nOut13_48), .ScanIn(nScanOut945), .ScanOut(nScanOut944), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_945 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_49), .NorthIn(nOut14_48), .SouthIn(nOut14_50), .EastIn(nOut15_49), .WestIn(nOut13_49), .ScanIn(nScanOut946), .ScanOut(nScanOut945), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_946 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_50), .NorthIn(nOut14_49), .SouthIn(nOut14_51), .EastIn(nOut15_50), .WestIn(nOut13_50), .ScanIn(nScanOut947), .ScanOut(nScanOut946), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_947 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_51), .NorthIn(nOut14_50), .SouthIn(nOut14_52), .EastIn(nOut15_51), .WestIn(nOut13_51), .ScanIn(nScanOut948), .ScanOut(nScanOut947), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_948 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_52), .NorthIn(nOut14_51), .SouthIn(nOut14_53), .EastIn(nOut15_52), .WestIn(nOut13_52), .ScanIn(nScanOut949), .ScanOut(nScanOut948), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_949 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_53), .NorthIn(nOut14_52), .SouthIn(nOut14_54), .EastIn(nOut15_53), .WestIn(nOut13_53), .ScanIn(nScanOut950), .ScanOut(nScanOut949), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_950 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_54), .NorthIn(nOut14_53), .SouthIn(nOut14_55), .EastIn(nOut15_54), .WestIn(nOut13_54), .ScanIn(nScanOut951), .ScanOut(nScanOut950), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_951 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_55), .NorthIn(nOut14_54), .SouthIn(nOut14_56), .EastIn(nOut15_55), .WestIn(nOut13_55), .ScanIn(nScanOut952), .ScanOut(nScanOut951), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_952 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_56), .NorthIn(nOut14_55), .SouthIn(nOut14_57), .EastIn(nOut15_56), .WestIn(nOut13_56), .ScanIn(nScanOut953), .ScanOut(nScanOut952), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_953 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_57), .NorthIn(nOut14_56), .SouthIn(nOut14_58), .EastIn(nOut15_57), .WestIn(nOut13_57), .ScanIn(nScanOut954), .ScanOut(nScanOut953), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_954 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_58), .NorthIn(nOut14_57), .SouthIn(nOut14_59), .EastIn(nOut15_58), .WestIn(nOut13_58), .ScanIn(nScanOut955), .ScanOut(nScanOut954), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_955 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_59), .NorthIn(nOut14_58), .SouthIn(nOut14_60), .EastIn(nOut15_59), .WestIn(nOut13_59), .ScanIn(nScanOut956), .ScanOut(nScanOut955), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_956 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_60), .NorthIn(nOut14_59), .SouthIn(nOut14_61), .EastIn(nOut15_60), .WestIn(nOut13_60), .ScanIn(nScanOut957), .ScanOut(nScanOut956), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_957 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_61), .NorthIn(nOut14_60), .SouthIn(nOut14_62), .EastIn(nOut15_61), .WestIn(nOut13_61), .ScanIn(nScanOut958), .ScanOut(nScanOut957), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_958 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_62), .NorthIn(nOut14_61), .SouthIn(nOut14_63), .EastIn(nOut15_62), .WestIn(nOut13_62), .ScanIn(nScanOut959), .ScanOut(nScanOut958), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_959 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut14_63), .ScanIn(nScanOut960), .ScanOut(nScanOut959), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_960 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_0), .ScanIn(nScanOut961), .ScanOut(nScanOut960), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_961 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_1), .NorthIn(nOut15_0), .SouthIn(nOut15_2), .EastIn(nOut16_1), .WestIn(nOut14_1), .ScanIn(nScanOut962), .ScanOut(nScanOut961), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_962 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_2), .NorthIn(nOut15_1), .SouthIn(nOut15_3), .EastIn(nOut16_2), .WestIn(nOut14_2), .ScanIn(nScanOut963), .ScanOut(nScanOut962), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_963 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_3), .NorthIn(nOut15_2), .SouthIn(nOut15_4), .EastIn(nOut16_3), .WestIn(nOut14_3), .ScanIn(nScanOut964), .ScanOut(nScanOut963), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_964 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_4), .NorthIn(nOut15_3), .SouthIn(nOut15_5), .EastIn(nOut16_4), .WestIn(nOut14_4), .ScanIn(nScanOut965), .ScanOut(nScanOut964), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_965 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_5), .NorthIn(nOut15_4), .SouthIn(nOut15_6), .EastIn(nOut16_5), .WestIn(nOut14_5), .ScanIn(nScanOut966), .ScanOut(nScanOut965), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_966 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_6), .NorthIn(nOut15_5), .SouthIn(nOut15_7), .EastIn(nOut16_6), .WestIn(nOut14_6), .ScanIn(nScanOut967), .ScanOut(nScanOut966), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_967 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_7), .NorthIn(nOut15_6), .SouthIn(nOut15_8), .EastIn(nOut16_7), .WestIn(nOut14_7), .ScanIn(nScanOut968), .ScanOut(nScanOut967), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_968 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_8), .NorthIn(nOut15_7), .SouthIn(nOut15_9), .EastIn(nOut16_8), .WestIn(nOut14_8), .ScanIn(nScanOut969), .ScanOut(nScanOut968), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_969 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_9), .NorthIn(nOut15_8), .SouthIn(nOut15_10), .EastIn(nOut16_9), .WestIn(nOut14_9), .ScanIn(nScanOut970), .ScanOut(nScanOut969), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_970 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_10), .NorthIn(nOut15_9), .SouthIn(nOut15_11), .EastIn(nOut16_10), .WestIn(nOut14_10), .ScanIn(nScanOut971), .ScanOut(nScanOut970), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_971 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_11), .NorthIn(nOut15_10), .SouthIn(nOut15_12), .EastIn(nOut16_11), .WestIn(nOut14_11), .ScanIn(nScanOut972), .ScanOut(nScanOut971), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_972 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_12), .NorthIn(nOut15_11), .SouthIn(nOut15_13), .EastIn(nOut16_12), .WestIn(nOut14_12), .ScanIn(nScanOut973), .ScanOut(nScanOut972), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_973 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_13), .NorthIn(nOut15_12), .SouthIn(nOut15_14), .EastIn(nOut16_13), .WestIn(nOut14_13), .ScanIn(nScanOut974), .ScanOut(nScanOut973), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_974 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_14), .NorthIn(nOut15_13), .SouthIn(nOut15_15), .EastIn(nOut16_14), .WestIn(nOut14_14), .ScanIn(nScanOut975), .ScanOut(nScanOut974), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_975 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_15), .NorthIn(nOut15_14), .SouthIn(nOut15_16), .EastIn(nOut16_15), .WestIn(nOut14_15), .ScanIn(nScanOut976), .ScanOut(nScanOut975), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_976 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_16), .NorthIn(nOut15_15), .SouthIn(nOut15_17), .EastIn(nOut16_16), .WestIn(nOut14_16), .ScanIn(nScanOut977), .ScanOut(nScanOut976), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_977 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_17), .NorthIn(nOut15_16), .SouthIn(nOut15_18), .EastIn(nOut16_17), .WestIn(nOut14_17), .ScanIn(nScanOut978), .ScanOut(nScanOut977), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_978 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_18), .NorthIn(nOut15_17), .SouthIn(nOut15_19), .EastIn(nOut16_18), .WestIn(nOut14_18), .ScanIn(nScanOut979), .ScanOut(nScanOut978), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_979 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_19), .NorthIn(nOut15_18), .SouthIn(nOut15_20), .EastIn(nOut16_19), .WestIn(nOut14_19), .ScanIn(nScanOut980), .ScanOut(nScanOut979), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_980 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_20), .NorthIn(nOut15_19), .SouthIn(nOut15_21), .EastIn(nOut16_20), .WestIn(nOut14_20), .ScanIn(nScanOut981), .ScanOut(nScanOut980), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_981 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_21), .NorthIn(nOut15_20), .SouthIn(nOut15_22), .EastIn(nOut16_21), .WestIn(nOut14_21), .ScanIn(nScanOut982), .ScanOut(nScanOut981), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_982 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_22), .NorthIn(nOut15_21), .SouthIn(nOut15_23), .EastIn(nOut16_22), .WestIn(nOut14_22), .ScanIn(nScanOut983), .ScanOut(nScanOut982), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_983 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_23), .NorthIn(nOut15_22), .SouthIn(nOut15_24), .EastIn(nOut16_23), .WestIn(nOut14_23), .ScanIn(nScanOut984), .ScanOut(nScanOut983), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_984 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_24), .NorthIn(nOut15_23), .SouthIn(nOut15_25), .EastIn(nOut16_24), .WestIn(nOut14_24), .ScanIn(nScanOut985), .ScanOut(nScanOut984), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_985 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_25), .NorthIn(nOut15_24), .SouthIn(nOut15_26), .EastIn(nOut16_25), .WestIn(nOut14_25), .ScanIn(nScanOut986), .ScanOut(nScanOut985), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_986 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_26), .NorthIn(nOut15_25), .SouthIn(nOut15_27), .EastIn(nOut16_26), .WestIn(nOut14_26), .ScanIn(nScanOut987), .ScanOut(nScanOut986), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_987 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_27), .NorthIn(nOut15_26), .SouthIn(nOut15_28), .EastIn(nOut16_27), .WestIn(nOut14_27), .ScanIn(nScanOut988), .ScanOut(nScanOut987), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_988 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_28), .NorthIn(nOut15_27), .SouthIn(nOut15_29), .EastIn(nOut16_28), .WestIn(nOut14_28), .ScanIn(nScanOut989), .ScanOut(nScanOut988), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_989 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_29), .NorthIn(nOut15_28), .SouthIn(nOut15_30), .EastIn(nOut16_29), .WestIn(nOut14_29), .ScanIn(nScanOut990), .ScanOut(nScanOut989), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_990 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_30), .NorthIn(nOut15_29), .SouthIn(nOut15_31), .EastIn(nOut16_30), .WestIn(nOut14_30), .ScanIn(nScanOut991), .ScanOut(nScanOut990), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_991 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_31), .NorthIn(nOut15_30), .SouthIn(nOut15_32), .EastIn(nOut16_31), .WestIn(nOut14_31), .ScanIn(nScanOut992), .ScanOut(nScanOut991), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_992 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_32), .NorthIn(nOut15_31), .SouthIn(nOut15_33), .EastIn(nOut16_32), .WestIn(nOut14_32), .ScanIn(nScanOut993), .ScanOut(nScanOut992), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_993 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_33), .NorthIn(nOut15_32), .SouthIn(nOut15_34), .EastIn(nOut16_33), .WestIn(nOut14_33), .ScanIn(nScanOut994), .ScanOut(nScanOut993), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_994 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_34), .NorthIn(nOut15_33), .SouthIn(nOut15_35), .EastIn(nOut16_34), .WestIn(nOut14_34), .ScanIn(nScanOut995), .ScanOut(nScanOut994), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_995 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_35), .NorthIn(nOut15_34), .SouthIn(nOut15_36), .EastIn(nOut16_35), .WestIn(nOut14_35), .ScanIn(nScanOut996), .ScanOut(nScanOut995), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_996 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_36), .NorthIn(nOut15_35), .SouthIn(nOut15_37), .EastIn(nOut16_36), .WestIn(nOut14_36), .ScanIn(nScanOut997), .ScanOut(nScanOut996), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_997 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_37), .NorthIn(nOut15_36), .SouthIn(nOut15_38), .EastIn(nOut16_37), .WestIn(nOut14_37), .ScanIn(nScanOut998), .ScanOut(nScanOut997), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_998 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_38), .NorthIn(nOut15_37), .SouthIn(nOut15_39), .EastIn(nOut16_38), .WestIn(nOut14_38), .ScanIn(nScanOut999), .ScanOut(nScanOut998), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_999 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_39), .NorthIn(nOut15_38), .SouthIn(nOut15_40), .EastIn(nOut16_39), .WestIn(nOut14_39), .ScanIn(nScanOut1000), .ScanOut(nScanOut999), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1000 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_40), .NorthIn(nOut15_39), .SouthIn(nOut15_41), .EastIn(nOut16_40), .WestIn(nOut14_40), .ScanIn(nScanOut1001), .ScanOut(nScanOut1000), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1001 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_41), .NorthIn(nOut15_40), .SouthIn(nOut15_42), .EastIn(nOut16_41), .WestIn(nOut14_41), .ScanIn(nScanOut1002), .ScanOut(nScanOut1001), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1002 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_42), .NorthIn(nOut15_41), .SouthIn(nOut15_43), .EastIn(nOut16_42), .WestIn(nOut14_42), .ScanIn(nScanOut1003), .ScanOut(nScanOut1002), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1003 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_43), .NorthIn(nOut15_42), .SouthIn(nOut15_44), .EastIn(nOut16_43), .WestIn(nOut14_43), .ScanIn(nScanOut1004), .ScanOut(nScanOut1003), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1004 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_44), .NorthIn(nOut15_43), .SouthIn(nOut15_45), .EastIn(nOut16_44), .WestIn(nOut14_44), .ScanIn(nScanOut1005), .ScanOut(nScanOut1004), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1005 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_45), .NorthIn(nOut15_44), .SouthIn(nOut15_46), .EastIn(nOut16_45), .WestIn(nOut14_45), .ScanIn(nScanOut1006), .ScanOut(nScanOut1005), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1006 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_46), .NorthIn(nOut15_45), .SouthIn(nOut15_47), .EastIn(nOut16_46), .WestIn(nOut14_46), .ScanIn(nScanOut1007), .ScanOut(nScanOut1006), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1007 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_47), .NorthIn(nOut15_46), .SouthIn(nOut15_48), .EastIn(nOut16_47), .WestIn(nOut14_47), .ScanIn(nScanOut1008), .ScanOut(nScanOut1007), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1008 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_48), .NorthIn(nOut15_47), .SouthIn(nOut15_49), .EastIn(nOut16_48), .WestIn(nOut14_48), .ScanIn(nScanOut1009), .ScanOut(nScanOut1008), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1009 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_49), .NorthIn(nOut15_48), .SouthIn(nOut15_50), .EastIn(nOut16_49), .WestIn(nOut14_49), .ScanIn(nScanOut1010), .ScanOut(nScanOut1009), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1010 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_50), .NorthIn(nOut15_49), .SouthIn(nOut15_51), .EastIn(nOut16_50), .WestIn(nOut14_50), .ScanIn(nScanOut1011), .ScanOut(nScanOut1010), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1011 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_51), .NorthIn(nOut15_50), .SouthIn(nOut15_52), .EastIn(nOut16_51), .WestIn(nOut14_51), .ScanIn(nScanOut1012), .ScanOut(nScanOut1011), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1012 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_52), .NorthIn(nOut15_51), .SouthIn(nOut15_53), .EastIn(nOut16_52), .WestIn(nOut14_52), .ScanIn(nScanOut1013), .ScanOut(nScanOut1012), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1013 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_53), .NorthIn(nOut15_52), .SouthIn(nOut15_54), .EastIn(nOut16_53), .WestIn(nOut14_53), .ScanIn(nScanOut1014), .ScanOut(nScanOut1013), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1014 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_54), .NorthIn(nOut15_53), .SouthIn(nOut15_55), .EastIn(nOut16_54), .WestIn(nOut14_54), .ScanIn(nScanOut1015), .ScanOut(nScanOut1014), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1015 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_55), .NorthIn(nOut15_54), .SouthIn(nOut15_56), .EastIn(nOut16_55), .WestIn(nOut14_55), .ScanIn(nScanOut1016), .ScanOut(nScanOut1015), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1016 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_56), .NorthIn(nOut15_55), .SouthIn(nOut15_57), .EastIn(nOut16_56), .WestIn(nOut14_56), .ScanIn(nScanOut1017), .ScanOut(nScanOut1016), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1017 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_57), .NorthIn(nOut15_56), .SouthIn(nOut15_58), .EastIn(nOut16_57), .WestIn(nOut14_57), .ScanIn(nScanOut1018), .ScanOut(nScanOut1017), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1018 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_58), .NorthIn(nOut15_57), .SouthIn(nOut15_59), .EastIn(nOut16_58), .WestIn(nOut14_58), .ScanIn(nScanOut1019), .ScanOut(nScanOut1018), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1019 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_59), .NorthIn(nOut15_58), .SouthIn(nOut15_60), .EastIn(nOut16_59), .WestIn(nOut14_59), .ScanIn(nScanOut1020), .ScanOut(nScanOut1019), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1020 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_60), .NorthIn(nOut15_59), .SouthIn(nOut15_61), .EastIn(nOut16_60), .WestIn(nOut14_60), .ScanIn(nScanOut1021), .ScanOut(nScanOut1020), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1021 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_61), .NorthIn(nOut15_60), .SouthIn(nOut15_62), .EastIn(nOut16_61), .WestIn(nOut14_61), .ScanIn(nScanOut1022), .ScanOut(nScanOut1021), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1022 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut15_62), .NorthIn(nOut15_61), .SouthIn(nOut15_63), .EastIn(nOut16_62), .WestIn(nOut14_62), .ScanIn(nScanOut1023), .ScanOut(nScanOut1022), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1023 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_63), .ScanIn(nScanOut1024), .ScanOut(nScanOut1023), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1024 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut16_0), .ScanIn(nScanOut1025), .ScanOut(nScanOut1024), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1025 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_1), .NorthIn(nOut16_0), .SouthIn(nOut16_2), .EastIn(nOut17_1), .WestIn(nOut15_1), .ScanIn(nScanOut1026), .ScanOut(nScanOut1025), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1026 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_2), .NorthIn(nOut16_1), .SouthIn(nOut16_3), .EastIn(nOut17_2), .WestIn(nOut15_2), .ScanIn(nScanOut1027), .ScanOut(nScanOut1026), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1027 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_3), .NorthIn(nOut16_2), .SouthIn(nOut16_4), .EastIn(nOut17_3), .WestIn(nOut15_3), .ScanIn(nScanOut1028), .ScanOut(nScanOut1027), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1028 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_4), .NorthIn(nOut16_3), .SouthIn(nOut16_5), .EastIn(nOut17_4), .WestIn(nOut15_4), .ScanIn(nScanOut1029), .ScanOut(nScanOut1028), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1029 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_5), .NorthIn(nOut16_4), .SouthIn(nOut16_6), .EastIn(nOut17_5), .WestIn(nOut15_5), .ScanIn(nScanOut1030), .ScanOut(nScanOut1029), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1030 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_6), .NorthIn(nOut16_5), .SouthIn(nOut16_7), .EastIn(nOut17_6), .WestIn(nOut15_6), .ScanIn(nScanOut1031), .ScanOut(nScanOut1030), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1031 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_7), .NorthIn(nOut16_6), .SouthIn(nOut16_8), .EastIn(nOut17_7), .WestIn(nOut15_7), .ScanIn(nScanOut1032), .ScanOut(nScanOut1031), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1032 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_8), .NorthIn(nOut16_7), .SouthIn(nOut16_9), .EastIn(nOut17_8), .WestIn(nOut15_8), .ScanIn(nScanOut1033), .ScanOut(nScanOut1032), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1033 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_9), .NorthIn(nOut16_8), .SouthIn(nOut16_10), .EastIn(nOut17_9), .WestIn(nOut15_9), .ScanIn(nScanOut1034), .ScanOut(nScanOut1033), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1034 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_10), .NorthIn(nOut16_9), .SouthIn(nOut16_11), .EastIn(nOut17_10), .WestIn(nOut15_10), .ScanIn(nScanOut1035), .ScanOut(nScanOut1034), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1035 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_11), .NorthIn(nOut16_10), .SouthIn(nOut16_12), .EastIn(nOut17_11), .WestIn(nOut15_11), .ScanIn(nScanOut1036), .ScanOut(nScanOut1035), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1036 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_12), .NorthIn(nOut16_11), .SouthIn(nOut16_13), .EastIn(nOut17_12), .WestIn(nOut15_12), .ScanIn(nScanOut1037), .ScanOut(nScanOut1036), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1037 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_13), .NorthIn(nOut16_12), .SouthIn(nOut16_14), .EastIn(nOut17_13), .WestIn(nOut15_13), .ScanIn(nScanOut1038), .ScanOut(nScanOut1037), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1038 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_14), .NorthIn(nOut16_13), .SouthIn(nOut16_15), .EastIn(nOut17_14), .WestIn(nOut15_14), .ScanIn(nScanOut1039), .ScanOut(nScanOut1038), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1039 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_15), .NorthIn(nOut16_14), .SouthIn(nOut16_16), .EastIn(nOut17_15), .WestIn(nOut15_15), .ScanIn(nScanOut1040), .ScanOut(nScanOut1039), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1040 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_16), .NorthIn(nOut16_15), .SouthIn(nOut16_17), .EastIn(nOut17_16), .WestIn(nOut15_16), .ScanIn(nScanOut1041), .ScanOut(nScanOut1040), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1041 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_17), .NorthIn(nOut16_16), .SouthIn(nOut16_18), .EastIn(nOut17_17), .WestIn(nOut15_17), .ScanIn(nScanOut1042), .ScanOut(nScanOut1041), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1042 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_18), .NorthIn(nOut16_17), .SouthIn(nOut16_19), .EastIn(nOut17_18), .WestIn(nOut15_18), .ScanIn(nScanOut1043), .ScanOut(nScanOut1042), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1043 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_19), .NorthIn(nOut16_18), .SouthIn(nOut16_20), .EastIn(nOut17_19), .WestIn(nOut15_19), .ScanIn(nScanOut1044), .ScanOut(nScanOut1043), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1044 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_20), .NorthIn(nOut16_19), .SouthIn(nOut16_21), .EastIn(nOut17_20), .WestIn(nOut15_20), .ScanIn(nScanOut1045), .ScanOut(nScanOut1044), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1045 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_21), .NorthIn(nOut16_20), .SouthIn(nOut16_22), .EastIn(nOut17_21), .WestIn(nOut15_21), .ScanIn(nScanOut1046), .ScanOut(nScanOut1045), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1046 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_22), .NorthIn(nOut16_21), .SouthIn(nOut16_23), .EastIn(nOut17_22), .WestIn(nOut15_22), .ScanIn(nScanOut1047), .ScanOut(nScanOut1046), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1047 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_23), .NorthIn(nOut16_22), .SouthIn(nOut16_24), .EastIn(nOut17_23), .WestIn(nOut15_23), .ScanIn(nScanOut1048), .ScanOut(nScanOut1047), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1048 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_24), .NorthIn(nOut16_23), .SouthIn(nOut16_25), .EastIn(nOut17_24), .WestIn(nOut15_24), .ScanIn(nScanOut1049), .ScanOut(nScanOut1048), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1049 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_25), .NorthIn(nOut16_24), .SouthIn(nOut16_26), .EastIn(nOut17_25), .WestIn(nOut15_25), .ScanIn(nScanOut1050), .ScanOut(nScanOut1049), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1050 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_26), .NorthIn(nOut16_25), .SouthIn(nOut16_27), .EastIn(nOut17_26), .WestIn(nOut15_26), .ScanIn(nScanOut1051), .ScanOut(nScanOut1050), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1051 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_27), .NorthIn(nOut16_26), .SouthIn(nOut16_28), .EastIn(nOut17_27), .WestIn(nOut15_27), .ScanIn(nScanOut1052), .ScanOut(nScanOut1051), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1052 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_28), .NorthIn(nOut16_27), .SouthIn(nOut16_29), .EastIn(nOut17_28), .WestIn(nOut15_28), .ScanIn(nScanOut1053), .ScanOut(nScanOut1052), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1053 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_29), .NorthIn(nOut16_28), .SouthIn(nOut16_30), .EastIn(nOut17_29), .WestIn(nOut15_29), .ScanIn(nScanOut1054), .ScanOut(nScanOut1053), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1054 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_30), .NorthIn(nOut16_29), .SouthIn(nOut16_31), .EastIn(nOut17_30), .WestIn(nOut15_30), .ScanIn(nScanOut1055), .ScanOut(nScanOut1054), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1055 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_31), .NorthIn(nOut16_30), .SouthIn(nOut16_32), .EastIn(nOut17_31), .WestIn(nOut15_31), .ScanIn(nScanOut1056), .ScanOut(nScanOut1055), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1056 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_32), .NorthIn(nOut16_31), .SouthIn(nOut16_33), .EastIn(nOut17_32), .WestIn(nOut15_32), .ScanIn(nScanOut1057), .ScanOut(nScanOut1056), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1057 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_33), .NorthIn(nOut16_32), .SouthIn(nOut16_34), .EastIn(nOut17_33), .WestIn(nOut15_33), .ScanIn(nScanOut1058), .ScanOut(nScanOut1057), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1058 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_34), .NorthIn(nOut16_33), .SouthIn(nOut16_35), .EastIn(nOut17_34), .WestIn(nOut15_34), .ScanIn(nScanOut1059), .ScanOut(nScanOut1058), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1059 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_35), .NorthIn(nOut16_34), .SouthIn(nOut16_36), .EastIn(nOut17_35), .WestIn(nOut15_35), .ScanIn(nScanOut1060), .ScanOut(nScanOut1059), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1060 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_36), .NorthIn(nOut16_35), .SouthIn(nOut16_37), .EastIn(nOut17_36), .WestIn(nOut15_36), .ScanIn(nScanOut1061), .ScanOut(nScanOut1060), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1061 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_37), .NorthIn(nOut16_36), .SouthIn(nOut16_38), .EastIn(nOut17_37), .WestIn(nOut15_37), .ScanIn(nScanOut1062), .ScanOut(nScanOut1061), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1062 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_38), .NorthIn(nOut16_37), .SouthIn(nOut16_39), .EastIn(nOut17_38), .WestIn(nOut15_38), .ScanIn(nScanOut1063), .ScanOut(nScanOut1062), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1063 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_39), .NorthIn(nOut16_38), .SouthIn(nOut16_40), .EastIn(nOut17_39), .WestIn(nOut15_39), .ScanIn(nScanOut1064), .ScanOut(nScanOut1063), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1064 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_40), .NorthIn(nOut16_39), .SouthIn(nOut16_41), .EastIn(nOut17_40), .WestIn(nOut15_40), .ScanIn(nScanOut1065), .ScanOut(nScanOut1064), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1065 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_41), .NorthIn(nOut16_40), .SouthIn(nOut16_42), .EastIn(nOut17_41), .WestIn(nOut15_41), .ScanIn(nScanOut1066), .ScanOut(nScanOut1065), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1066 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_42), .NorthIn(nOut16_41), .SouthIn(nOut16_43), .EastIn(nOut17_42), .WestIn(nOut15_42), .ScanIn(nScanOut1067), .ScanOut(nScanOut1066), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1067 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_43), .NorthIn(nOut16_42), .SouthIn(nOut16_44), .EastIn(nOut17_43), .WestIn(nOut15_43), .ScanIn(nScanOut1068), .ScanOut(nScanOut1067), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1068 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_44), .NorthIn(nOut16_43), .SouthIn(nOut16_45), .EastIn(nOut17_44), .WestIn(nOut15_44), .ScanIn(nScanOut1069), .ScanOut(nScanOut1068), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1069 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_45), .NorthIn(nOut16_44), .SouthIn(nOut16_46), .EastIn(nOut17_45), .WestIn(nOut15_45), .ScanIn(nScanOut1070), .ScanOut(nScanOut1069), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1070 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_46), .NorthIn(nOut16_45), .SouthIn(nOut16_47), .EastIn(nOut17_46), .WestIn(nOut15_46), .ScanIn(nScanOut1071), .ScanOut(nScanOut1070), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1071 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_47), .NorthIn(nOut16_46), .SouthIn(nOut16_48), .EastIn(nOut17_47), .WestIn(nOut15_47), .ScanIn(nScanOut1072), .ScanOut(nScanOut1071), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1072 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_48), .NorthIn(nOut16_47), .SouthIn(nOut16_49), .EastIn(nOut17_48), .WestIn(nOut15_48), .ScanIn(nScanOut1073), .ScanOut(nScanOut1072), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1073 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_49), .NorthIn(nOut16_48), .SouthIn(nOut16_50), .EastIn(nOut17_49), .WestIn(nOut15_49), .ScanIn(nScanOut1074), .ScanOut(nScanOut1073), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1074 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_50), .NorthIn(nOut16_49), .SouthIn(nOut16_51), .EastIn(nOut17_50), .WestIn(nOut15_50), .ScanIn(nScanOut1075), .ScanOut(nScanOut1074), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1075 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_51), .NorthIn(nOut16_50), .SouthIn(nOut16_52), .EastIn(nOut17_51), .WestIn(nOut15_51), .ScanIn(nScanOut1076), .ScanOut(nScanOut1075), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1076 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_52), .NorthIn(nOut16_51), .SouthIn(nOut16_53), .EastIn(nOut17_52), .WestIn(nOut15_52), .ScanIn(nScanOut1077), .ScanOut(nScanOut1076), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1077 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_53), .NorthIn(nOut16_52), .SouthIn(nOut16_54), .EastIn(nOut17_53), .WestIn(nOut15_53), .ScanIn(nScanOut1078), .ScanOut(nScanOut1077), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1078 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_54), .NorthIn(nOut16_53), .SouthIn(nOut16_55), .EastIn(nOut17_54), .WestIn(nOut15_54), .ScanIn(nScanOut1079), .ScanOut(nScanOut1078), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1079 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_55), .NorthIn(nOut16_54), .SouthIn(nOut16_56), .EastIn(nOut17_55), .WestIn(nOut15_55), .ScanIn(nScanOut1080), .ScanOut(nScanOut1079), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1080 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_56), .NorthIn(nOut16_55), .SouthIn(nOut16_57), .EastIn(nOut17_56), .WestIn(nOut15_56), .ScanIn(nScanOut1081), .ScanOut(nScanOut1080), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1081 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_57), .NorthIn(nOut16_56), .SouthIn(nOut16_58), .EastIn(nOut17_57), .WestIn(nOut15_57), .ScanIn(nScanOut1082), .ScanOut(nScanOut1081), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1082 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_58), .NorthIn(nOut16_57), .SouthIn(nOut16_59), .EastIn(nOut17_58), .WestIn(nOut15_58), .ScanIn(nScanOut1083), .ScanOut(nScanOut1082), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1083 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_59), .NorthIn(nOut16_58), .SouthIn(nOut16_60), .EastIn(nOut17_59), .WestIn(nOut15_59), .ScanIn(nScanOut1084), .ScanOut(nScanOut1083), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1084 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_60), .NorthIn(nOut16_59), .SouthIn(nOut16_61), .EastIn(nOut17_60), .WestIn(nOut15_60), .ScanIn(nScanOut1085), .ScanOut(nScanOut1084), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1085 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_61), .NorthIn(nOut16_60), .SouthIn(nOut16_62), .EastIn(nOut17_61), .WestIn(nOut15_61), .ScanIn(nScanOut1086), .ScanOut(nScanOut1085), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1086 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut16_62), .NorthIn(nOut16_61), .SouthIn(nOut16_63), .EastIn(nOut17_62), .WestIn(nOut15_62), .ScanIn(nScanOut1087), .ScanOut(nScanOut1086), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1087 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut16_63), .ScanIn(nScanOut1088), .ScanOut(nScanOut1087), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1088 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut17_0), .ScanIn(nScanOut1089), .ScanOut(nScanOut1088), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1089 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_1), .NorthIn(nOut17_0), .SouthIn(nOut17_2), .EastIn(nOut18_1), .WestIn(nOut16_1), .ScanIn(nScanOut1090), .ScanOut(nScanOut1089), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1090 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_2), .NorthIn(nOut17_1), .SouthIn(nOut17_3), .EastIn(nOut18_2), .WestIn(nOut16_2), .ScanIn(nScanOut1091), .ScanOut(nScanOut1090), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1091 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_3), .NorthIn(nOut17_2), .SouthIn(nOut17_4), .EastIn(nOut18_3), .WestIn(nOut16_3), .ScanIn(nScanOut1092), .ScanOut(nScanOut1091), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1092 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_4), .NorthIn(nOut17_3), .SouthIn(nOut17_5), .EastIn(nOut18_4), .WestIn(nOut16_4), .ScanIn(nScanOut1093), .ScanOut(nScanOut1092), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1093 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_5), .NorthIn(nOut17_4), .SouthIn(nOut17_6), .EastIn(nOut18_5), .WestIn(nOut16_5), .ScanIn(nScanOut1094), .ScanOut(nScanOut1093), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1094 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_6), .NorthIn(nOut17_5), .SouthIn(nOut17_7), .EastIn(nOut18_6), .WestIn(nOut16_6), .ScanIn(nScanOut1095), .ScanOut(nScanOut1094), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1095 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_7), .NorthIn(nOut17_6), .SouthIn(nOut17_8), .EastIn(nOut18_7), .WestIn(nOut16_7), .ScanIn(nScanOut1096), .ScanOut(nScanOut1095), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1096 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_8), .NorthIn(nOut17_7), .SouthIn(nOut17_9), .EastIn(nOut18_8), .WestIn(nOut16_8), .ScanIn(nScanOut1097), .ScanOut(nScanOut1096), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1097 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_9), .NorthIn(nOut17_8), .SouthIn(nOut17_10), .EastIn(nOut18_9), .WestIn(nOut16_9), .ScanIn(nScanOut1098), .ScanOut(nScanOut1097), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1098 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_10), .NorthIn(nOut17_9), .SouthIn(nOut17_11), .EastIn(nOut18_10), .WestIn(nOut16_10), .ScanIn(nScanOut1099), .ScanOut(nScanOut1098), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1099 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_11), .NorthIn(nOut17_10), .SouthIn(nOut17_12), .EastIn(nOut18_11), .WestIn(nOut16_11), .ScanIn(nScanOut1100), .ScanOut(nScanOut1099), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_12), .NorthIn(nOut17_11), .SouthIn(nOut17_13), .EastIn(nOut18_12), .WestIn(nOut16_12), .ScanIn(nScanOut1101), .ScanOut(nScanOut1100), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_13), .NorthIn(nOut17_12), .SouthIn(nOut17_14), .EastIn(nOut18_13), .WestIn(nOut16_13), .ScanIn(nScanOut1102), .ScanOut(nScanOut1101), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_14), .NorthIn(nOut17_13), .SouthIn(nOut17_15), .EastIn(nOut18_14), .WestIn(nOut16_14), .ScanIn(nScanOut1103), .ScanOut(nScanOut1102), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_15), .NorthIn(nOut17_14), .SouthIn(nOut17_16), .EastIn(nOut18_15), .WestIn(nOut16_15), .ScanIn(nScanOut1104), .ScanOut(nScanOut1103), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_16), .NorthIn(nOut17_15), .SouthIn(nOut17_17), .EastIn(nOut18_16), .WestIn(nOut16_16), .ScanIn(nScanOut1105), .ScanOut(nScanOut1104), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_17), .NorthIn(nOut17_16), .SouthIn(nOut17_18), .EastIn(nOut18_17), .WestIn(nOut16_17), .ScanIn(nScanOut1106), .ScanOut(nScanOut1105), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_18), .NorthIn(nOut17_17), .SouthIn(nOut17_19), .EastIn(nOut18_18), .WestIn(nOut16_18), .ScanIn(nScanOut1107), .ScanOut(nScanOut1106), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_19), .NorthIn(nOut17_18), .SouthIn(nOut17_20), .EastIn(nOut18_19), .WestIn(nOut16_19), .ScanIn(nScanOut1108), .ScanOut(nScanOut1107), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_20), .NorthIn(nOut17_19), .SouthIn(nOut17_21), .EastIn(nOut18_20), .WestIn(nOut16_20), .ScanIn(nScanOut1109), .ScanOut(nScanOut1108), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_21), .NorthIn(nOut17_20), .SouthIn(nOut17_22), .EastIn(nOut18_21), .WestIn(nOut16_21), .ScanIn(nScanOut1110), .ScanOut(nScanOut1109), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_22), .NorthIn(nOut17_21), .SouthIn(nOut17_23), .EastIn(nOut18_22), .WestIn(nOut16_22), .ScanIn(nScanOut1111), .ScanOut(nScanOut1110), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_23), .NorthIn(nOut17_22), .SouthIn(nOut17_24), .EastIn(nOut18_23), .WestIn(nOut16_23), .ScanIn(nScanOut1112), .ScanOut(nScanOut1111), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_24), .NorthIn(nOut17_23), .SouthIn(nOut17_25), .EastIn(nOut18_24), .WestIn(nOut16_24), .ScanIn(nScanOut1113), .ScanOut(nScanOut1112), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_25), .NorthIn(nOut17_24), .SouthIn(nOut17_26), .EastIn(nOut18_25), .WestIn(nOut16_25), .ScanIn(nScanOut1114), .ScanOut(nScanOut1113), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_26), .NorthIn(nOut17_25), .SouthIn(nOut17_27), .EastIn(nOut18_26), .WestIn(nOut16_26), .ScanIn(nScanOut1115), .ScanOut(nScanOut1114), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_27), .NorthIn(nOut17_26), .SouthIn(nOut17_28), .EastIn(nOut18_27), .WestIn(nOut16_27), .ScanIn(nScanOut1116), .ScanOut(nScanOut1115), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_28), .NorthIn(nOut17_27), .SouthIn(nOut17_29), .EastIn(nOut18_28), .WestIn(nOut16_28), .ScanIn(nScanOut1117), .ScanOut(nScanOut1116), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_29), .NorthIn(nOut17_28), .SouthIn(nOut17_30), .EastIn(nOut18_29), .WestIn(nOut16_29), .ScanIn(nScanOut1118), .ScanOut(nScanOut1117), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_30), .NorthIn(nOut17_29), .SouthIn(nOut17_31), .EastIn(nOut18_30), .WestIn(nOut16_30), .ScanIn(nScanOut1119), .ScanOut(nScanOut1118), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_31), .NorthIn(nOut17_30), .SouthIn(nOut17_32), .EastIn(nOut18_31), .WestIn(nOut16_31), .ScanIn(nScanOut1120), .ScanOut(nScanOut1119), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_32), .NorthIn(nOut17_31), .SouthIn(nOut17_33), .EastIn(nOut18_32), .WestIn(nOut16_32), .ScanIn(nScanOut1121), .ScanOut(nScanOut1120), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_33), .NorthIn(nOut17_32), .SouthIn(nOut17_34), .EastIn(nOut18_33), .WestIn(nOut16_33), .ScanIn(nScanOut1122), .ScanOut(nScanOut1121), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_34), .NorthIn(nOut17_33), .SouthIn(nOut17_35), .EastIn(nOut18_34), .WestIn(nOut16_34), .ScanIn(nScanOut1123), .ScanOut(nScanOut1122), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_35), .NorthIn(nOut17_34), .SouthIn(nOut17_36), .EastIn(nOut18_35), .WestIn(nOut16_35), .ScanIn(nScanOut1124), .ScanOut(nScanOut1123), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_36), .NorthIn(nOut17_35), .SouthIn(nOut17_37), .EastIn(nOut18_36), .WestIn(nOut16_36), .ScanIn(nScanOut1125), .ScanOut(nScanOut1124), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_37), .NorthIn(nOut17_36), .SouthIn(nOut17_38), .EastIn(nOut18_37), .WestIn(nOut16_37), .ScanIn(nScanOut1126), .ScanOut(nScanOut1125), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_38), .NorthIn(nOut17_37), .SouthIn(nOut17_39), .EastIn(nOut18_38), .WestIn(nOut16_38), .ScanIn(nScanOut1127), .ScanOut(nScanOut1126), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_39), .NorthIn(nOut17_38), .SouthIn(nOut17_40), .EastIn(nOut18_39), .WestIn(nOut16_39), .ScanIn(nScanOut1128), .ScanOut(nScanOut1127), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_40), .NorthIn(nOut17_39), .SouthIn(nOut17_41), .EastIn(nOut18_40), .WestIn(nOut16_40), .ScanIn(nScanOut1129), .ScanOut(nScanOut1128), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_41), .NorthIn(nOut17_40), .SouthIn(nOut17_42), .EastIn(nOut18_41), .WestIn(nOut16_41), .ScanIn(nScanOut1130), .ScanOut(nScanOut1129), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_42), .NorthIn(nOut17_41), .SouthIn(nOut17_43), .EastIn(nOut18_42), .WestIn(nOut16_42), .ScanIn(nScanOut1131), .ScanOut(nScanOut1130), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_43), .NorthIn(nOut17_42), .SouthIn(nOut17_44), .EastIn(nOut18_43), .WestIn(nOut16_43), .ScanIn(nScanOut1132), .ScanOut(nScanOut1131), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_44), .NorthIn(nOut17_43), .SouthIn(nOut17_45), .EastIn(nOut18_44), .WestIn(nOut16_44), .ScanIn(nScanOut1133), .ScanOut(nScanOut1132), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_45), .NorthIn(nOut17_44), .SouthIn(nOut17_46), .EastIn(nOut18_45), .WestIn(nOut16_45), .ScanIn(nScanOut1134), .ScanOut(nScanOut1133), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_46), .NorthIn(nOut17_45), .SouthIn(nOut17_47), .EastIn(nOut18_46), .WestIn(nOut16_46), .ScanIn(nScanOut1135), .ScanOut(nScanOut1134), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_47), .NorthIn(nOut17_46), .SouthIn(nOut17_48), .EastIn(nOut18_47), .WestIn(nOut16_47), .ScanIn(nScanOut1136), .ScanOut(nScanOut1135), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_48), .NorthIn(nOut17_47), .SouthIn(nOut17_49), .EastIn(nOut18_48), .WestIn(nOut16_48), .ScanIn(nScanOut1137), .ScanOut(nScanOut1136), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_49), .NorthIn(nOut17_48), .SouthIn(nOut17_50), .EastIn(nOut18_49), .WestIn(nOut16_49), .ScanIn(nScanOut1138), .ScanOut(nScanOut1137), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_50), .NorthIn(nOut17_49), .SouthIn(nOut17_51), .EastIn(nOut18_50), .WestIn(nOut16_50), .ScanIn(nScanOut1139), .ScanOut(nScanOut1138), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_51), .NorthIn(nOut17_50), .SouthIn(nOut17_52), .EastIn(nOut18_51), .WestIn(nOut16_51), .ScanIn(nScanOut1140), .ScanOut(nScanOut1139), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_52), .NorthIn(nOut17_51), .SouthIn(nOut17_53), .EastIn(nOut18_52), .WestIn(nOut16_52), .ScanIn(nScanOut1141), .ScanOut(nScanOut1140), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_53), .NorthIn(nOut17_52), .SouthIn(nOut17_54), .EastIn(nOut18_53), .WestIn(nOut16_53), .ScanIn(nScanOut1142), .ScanOut(nScanOut1141), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_54), .NorthIn(nOut17_53), .SouthIn(nOut17_55), .EastIn(nOut18_54), .WestIn(nOut16_54), .ScanIn(nScanOut1143), .ScanOut(nScanOut1142), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_55), .NorthIn(nOut17_54), .SouthIn(nOut17_56), .EastIn(nOut18_55), .WestIn(nOut16_55), .ScanIn(nScanOut1144), .ScanOut(nScanOut1143), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_56), .NorthIn(nOut17_55), .SouthIn(nOut17_57), .EastIn(nOut18_56), .WestIn(nOut16_56), .ScanIn(nScanOut1145), .ScanOut(nScanOut1144), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_57), .NorthIn(nOut17_56), .SouthIn(nOut17_58), .EastIn(nOut18_57), .WestIn(nOut16_57), .ScanIn(nScanOut1146), .ScanOut(nScanOut1145), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_58), .NorthIn(nOut17_57), .SouthIn(nOut17_59), .EastIn(nOut18_58), .WestIn(nOut16_58), .ScanIn(nScanOut1147), .ScanOut(nScanOut1146), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_59), .NorthIn(nOut17_58), .SouthIn(nOut17_60), .EastIn(nOut18_59), .WestIn(nOut16_59), .ScanIn(nScanOut1148), .ScanOut(nScanOut1147), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_60), .NorthIn(nOut17_59), .SouthIn(nOut17_61), .EastIn(nOut18_60), .WestIn(nOut16_60), .ScanIn(nScanOut1149), .ScanOut(nScanOut1148), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_61), .NorthIn(nOut17_60), .SouthIn(nOut17_62), .EastIn(nOut18_61), .WestIn(nOut16_61), .ScanIn(nScanOut1150), .ScanOut(nScanOut1149), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut17_62), .NorthIn(nOut17_61), .SouthIn(nOut17_63), .EastIn(nOut18_62), .WestIn(nOut16_62), .ScanIn(nScanOut1151), .ScanOut(nScanOut1150), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut17_63), .ScanIn(nScanOut1152), .ScanOut(nScanOut1151), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut18_0), .ScanIn(nScanOut1153), .ScanOut(nScanOut1152), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_1), .NorthIn(nOut18_0), .SouthIn(nOut18_2), .EastIn(nOut19_1), .WestIn(nOut17_1), .ScanIn(nScanOut1154), .ScanOut(nScanOut1153), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_2), .NorthIn(nOut18_1), .SouthIn(nOut18_3), .EastIn(nOut19_2), .WestIn(nOut17_2), .ScanIn(nScanOut1155), .ScanOut(nScanOut1154), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_3), .NorthIn(nOut18_2), .SouthIn(nOut18_4), .EastIn(nOut19_3), .WestIn(nOut17_3), .ScanIn(nScanOut1156), .ScanOut(nScanOut1155), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_4), .NorthIn(nOut18_3), .SouthIn(nOut18_5), .EastIn(nOut19_4), .WestIn(nOut17_4), .ScanIn(nScanOut1157), .ScanOut(nScanOut1156), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_5), .NorthIn(nOut18_4), .SouthIn(nOut18_6), .EastIn(nOut19_5), .WestIn(nOut17_5), .ScanIn(nScanOut1158), .ScanOut(nScanOut1157), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_6), .NorthIn(nOut18_5), .SouthIn(nOut18_7), .EastIn(nOut19_6), .WestIn(nOut17_6), .ScanIn(nScanOut1159), .ScanOut(nScanOut1158), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_7), .NorthIn(nOut18_6), .SouthIn(nOut18_8), .EastIn(nOut19_7), .WestIn(nOut17_7), .ScanIn(nScanOut1160), .ScanOut(nScanOut1159), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_8), .NorthIn(nOut18_7), .SouthIn(nOut18_9), .EastIn(nOut19_8), .WestIn(nOut17_8), .ScanIn(nScanOut1161), .ScanOut(nScanOut1160), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_9), .NorthIn(nOut18_8), .SouthIn(nOut18_10), .EastIn(nOut19_9), .WestIn(nOut17_9), .ScanIn(nScanOut1162), .ScanOut(nScanOut1161), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_10), .NorthIn(nOut18_9), .SouthIn(nOut18_11), .EastIn(nOut19_10), .WestIn(nOut17_10), .ScanIn(nScanOut1163), .ScanOut(nScanOut1162), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_11), .NorthIn(nOut18_10), .SouthIn(nOut18_12), .EastIn(nOut19_11), .WestIn(nOut17_11), .ScanIn(nScanOut1164), .ScanOut(nScanOut1163), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_12), .NorthIn(nOut18_11), .SouthIn(nOut18_13), .EastIn(nOut19_12), .WestIn(nOut17_12), .ScanIn(nScanOut1165), .ScanOut(nScanOut1164), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_13), .NorthIn(nOut18_12), .SouthIn(nOut18_14), .EastIn(nOut19_13), .WestIn(nOut17_13), .ScanIn(nScanOut1166), .ScanOut(nScanOut1165), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_14), .NorthIn(nOut18_13), .SouthIn(nOut18_15), .EastIn(nOut19_14), .WestIn(nOut17_14), .ScanIn(nScanOut1167), .ScanOut(nScanOut1166), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_15), .NorthIn(nOut18_14), .SouthIn(nOut18_16), .EastIn(nOut19_15), .WestIn(nOut17_15), .ScanIn(nScanOut1168), .ScanOut(nScanOut1167), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_16), .NorthIn(nOut18_15), .SouthIn(nOut18_17), .EastIn(nOut19_16), .WestIn(nOut17_16), .ScanIn(nScanOut1169), .ScanOut(nScanOut1168), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_17), .NorthIn(nOut18_16), .SouthIn(nOut18_18), .EastIn(nOut19_17), .WestIn(nOut17_17), .ScanIn(nScanOut1170), .ScanOut(nScanOut1169), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_18), .NorthIn(nOut18_17), .SouthIn(nOut18_19), .EastIn(nOut19_18), .WestIn(nOut17_18), .ScanIn(nScanOut1171), .ScanOut(nScanOut1170), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_19), .NorthIn(nOut18_18), .SouthIn(nOut18_20), .EastIn(nOut19_19), .WestIn(nOut17_19), .ScanIn(nScanOut1172), .ScanOut(nScanOut1171), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_20), .NorthIn(nOut18_19), .SouthIn(nOut18_21), .EastIn(nOut19_20), .WestIn(nOut17_20), .ScanIn(nScanOut1173), .ScanOut(nScanOut1172), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_21), .NorthIn(nOut18_20), .SouthIn(nOut18_22), .EastIn(nOut19_21), .WestIn(nOut17_21), .ScanIn(nScanOut1174), .ScanOut(nScanOut1173), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_22), .NorthIn(nOut18_21), .SouthIn(nOut18_23), .EastIn(nOut19_22), .WestIn(nOut17_22), .ScanIn(nScanOut1175), .ScanOut(nScanOut1174), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_23), .NorthIn(nOut18_22), .SouthIn(nOut18_24), .EastIn(nOut19_23), .WestIn(nOut17_23), .ScanIn(nScanOut1176), .ScanOut(nScanOut1175), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_24), .NorthIn(nOut18_23), .SouthIn(nOut18_25), .EastIn(nOut19_24), .WestIn(nOut17_24), .ScanIn(nScanOut1177), .ScanOut(nScanOut1176), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_25), .NorthIn(nOut18_24), .SouthIn(nOut18_26), .EastIn(nOut19_25), .WestIn(nOut17_25), .ScanIn(nScanOut1178), .ScanOut(nScanOut1177), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_26), .NorthIn(nOut18_25), .SouthIn(nOut18_27), .EastIn(nOut19_26), .WestIn(nOut17_26), .ScanIn(nScanOut1179), .ScanOut(nScanOut1178), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_27), .NorthIn(nOut18_26), .SouthIn(nOut18_28), .EastIn(nOut19_27), .WestIn(nOut17_27), .ScanIn(nScanOut1180), .ScanOut(nScanOut1179), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_28), .NorthIn(nOut18_27), .SouthIn(nOut18_29), .EastIn(nOut19_28), .WestIn(nOut17_28), .ScanIn(nScanOut1181), .ScanOut(nScanOut1180), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_29), .NorthIn(nOut18_28), .SouthIn(nOut18_30), .EastIn(nOut19_29), .WestIn(nOut17_29), .ScanIn(nScanOut1182), .ScanOut(nScanOut1181), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_30), .NorthIn(nOut18_29), .SouthIn(nOut18_31), .EastIn(nOut19_30), .WestIn(nOut17_30), .ScanIn(nScanOut1183), .ScanOut(nScanOut1182), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_31), .NorthIn(nOut18_30), .SouthIn(nOut18_32), .EastIn(nOut19_31), .WestIn(nOut17_31), .ScanIn(nScanOut1184), .ScanOut(nScanOut1183), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_32), .NorthIn(nOut18_31), .SouthIn(nOut18_33), .EastIn(nOut19_32), .WestIn(nOut17_32), .ScanIn(nScanOut1185), .ScanOut(nScanOut1184), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_33), .NorthIn(nOut18_32), .SouthIn(nOut18_34), .EastIn(nOut19_33), .WestIn(nOut17_33), .ScanIn(nScanOut1186), .ScanOut(nScanOut1185), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_34), .NorthIn(nOut18_33), .SouthIn(nOut18_35), .EastIn(nOut19_34), .WestIn(nOut17_34), .ScanIn(nScanOut1187), .ScanOut(nScanOut1186), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_35), .NorthIn(nOut18_34), .SouthIn(nOut18_36), .EastIn(nOut19_35), .WestIn(nOut17_35), .ScanIn(nScanOut1188), .ScanOut(nScanOut1187), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_36), .NorthIn(nOut18_35), .SouthIn(nOut18_37), .EastIn(nOut19_36), .WestIn(nOut17_36), .ScanIn(nScanOut1189), .ScanOut(nScanOut1188), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_37), .NorthIn(nOut18_36), .SouthIn(nOut18_38), .EastIn(nOut19_37), .WestIn(nOut17_37), .ScanIn(nScanOut1190), .ScanOut(nScanOut1189), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_38), .NorthIn(nOut18_37), .SouthIn(nOut18_39), .EastIn(nOut19_38), .WestIn(nOut17_38), .ScanIn(nScanOut1191), .ScanOut(nScanOut1190), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_39), .NorthIn(nOut18_38), .SouthIn(nOut18_40), .EastIn(nOut19_39), .WestIn(nOut17_39), .ScanIn(nScanOut1192), .ScanOut(nScanOut1191), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_40), .NorthIn(nOut18_39), .SouthIn(nOut18_41), .EastIn(nOut19_40), .WestIn(nOut17_40), .ScanIn(nScanOut1193), .ScanOut(nScanOut1192), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_41), .NorthIn(nOut18_40), .SouthIn(nOut18_42), .EastIn(nOut19_41), .WestIn(nOut17_41), .ScanIn(nScanOut1194), .ScanOut(nScanOut1193), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_42), .NorthIn(nOut18_41), .SouthIn(nOut18_43), .EastIn(nOut19_42), .WestIn(nOut17_42), .ScanIn(nScanOut1195), .ScanOut(nScanOut1194), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_43), .NorthIn(nOut18_42), .SouthIn(nOut18_44), .EastIn(nOut19_43), .WestIn(nOut17_43), .ScanIn(nScanOut1196), .ScanOut(nScanOut1195), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_44), .NorthIn(nOut18_43), .SouthIn(nOut18_45), .EastIn(nOut19_44), .WestIn(nOut17_44), .ScanIn(nScanOut1197), .ScanOut(nScanOut1196), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_45), .NorthIn(nOut18_44), .SouthIn(nOut18_46), .EastIn(nOut19_45), .WestIn(nOut17_45), .ScanIn(nScanOut1198), .ScanOut(nScanOut1197), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_46), .NorthIn(nOut18_45), .SouthIn(nOut18_47), .EastIn(nOut19_46), .WestIn(nOut17_46), .ScanIn(nScanOut1199), .ScanOut(nScanOut1198), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_47), .NorthIn(nOut18_46), .SouthIn(nOut18_48), .EastIn(nOut19_47), .WestIn(nOut17_47), .ScanIn(nScanOut1200), .ScanOut(nScanOut1199), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_48), .NorthIn(nOut18_47), .SouthIn(nOut18_49), .EastIn(nOut19_48), .WestIn(nOut17_48), .ScanIn(nScanOut1201), .ScanOut(nScanOut1200), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_49), .NorthIn(nOut18_48), .SouthIn(nOut18_50), .EastIn(nOut19_49), .WestIn(nOut17_49), .ScanIn(nScanOut1202), .ScanOut(nScanOut1201), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_50), .NorthIn(nOut18_49), .SouthIn(nOut18_51), .EastIn(nOut19_50), .WestIn(nOut17_50), .ScanIn(nScanOut1203), .ScanOut(nScanOut1202), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_51), .NorthIn(nOut18_50), .SouthIn(nOut18_52), .EastIn(nOut19_51), .WestIn(nOut17_51), .ScanIn(nScanOut1204), .ScanOut(nScanOut1203), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_52), .NorthIn(nOut18_51), .SouthIn(nOut18_53), .EastIn(nOut19_52), .WestIn(nOut17_52), .ScanIn(nScanOut1205), .ScanOut(nScanOut1204), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_53), .NorthIn(nOut18_52), .SouthIn(nOut18_54), .EastIn(nOut19_53), .WestIn(nOut17_53), .ScanIn(nScanOut1206), .ScanOut(nScanOut1205), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_54), .NorthIn(nOut18_53), .SouthIn(nOut18_55), .EastIn(nOut19_54), .WestIn(nOut17_54), .ScanIn(nScanOut1207), .ScanOut(nScanOut1206), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_55), .NorthIn(nOut18_54), .SouthIn(nOut18_56), .EastIn(nOut19_55), .WestIn(nOut17_55), .ScanIn(nScanOut1208), .ScanOut(nScanOut1207), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_56), .NorthIn(nOut18_55), .SouthIn(nOut18_57), .EastIn(nOut19_56), .WestIn(nOut17_56), .ScanIn(nScanOut1209), .ScanOut(nScanOut1208), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_57), .NorthIn(nOut18_56), .SouthIn(nOut18_58), .EastIn(nOut19_57), .WestIn(nOut17_57), .ScanIn(nScanOut1210), .ScanOut(nScanOut1209), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_58), .NorthIn(nOut18_57), .SouthIn(nOut18_59), .EastIn(nOut19_58), .WestIn(nOut17_58), .ScanIn(nScanOut1211), .ScanOut(nScanOut1210), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_59), .NorthIn(nOut18_58), .SouthIn(nOut18_60), .EastIn(nOut19_59), .WestIn(nOut17_59), .ScanIn(nScanOut1212), .ScanOut(nScanOut1211), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_60), .NorthIn(nOut18_59), .SouthIn(nOut18_61), .EastIn(nOut19_60), .WestIn(nOut17_60), .ScanIn(nScanOut1213), .ScanOut(nScanOut1212), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_61), .NorthIn(nOut18_60), .SouthIn(nOut18_62), .EastIn(nOut19_61), .WestIn(nOut17_61), .ScanIn(nScanOut1214), .ScanOut(nScanOut1213), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut18_62), .NorthIn(nOut18_61), .SouthIn(nOut18_63), .EastIn(nOut19_62), .WestIn(nOut17_62), .ScanIn(nScanOut1215), .ScanOut(nScanOut1214), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut18_63), .ScanIn(nScanOut1216), .ScanOut(nScanOut1215), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut19_0), .ScanIn(nScanOut1217), .ScanOut(nScanOut1216), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_1), .NorthIn(nOut19_0), .SouthIn(nOut19_2), .EastIn(nOut20_1), .WestIn(nOut18_1), .ScanIn(nScanOut1218), .ScanOut(nScanOut1217), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_2), .NorthIn(nOut19_1), .SouthIn(nOut19_3), .EastIn(nOut20_2), .WestIn(nOut18_2), .ScanIn(nScanOut1219), .ScanOut(nScanOut1218), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_3), .NorthIn(nOut19_2), .SouthIn(nOut19_4), .EastIn(nOut20_3), .WestIn(nOut18_3), .ScanIn(nScanOut1220), .ScanOut(nScanOut1219), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_4), .NorthIn(nOut19_3), .SouthIn(nOut19_5), .EastIn(nOut20_4), .WestIn(nOut18_4), .ScanIn(nScanOut1221), .ScanOut(nScanOut1220), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_5), .NorthIn(nOut19_4), .SouthIn(nOut19_6), .EastIn(nOut20_5), .WestIn(nOut18_5), .ScanIn(nScanOut1222), .ScanOut(nScanOut1221), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_6), .NorthIn(nOut19_5), .SouthIn(nOut19_7), .EastIn(nOut20_6), .WestIn(nOut18_6), .ScanIn(nScanOut1223), .ScanOut(nScanOut1222), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_7), .NorthIn(nOut19_6), .SouthIn(nOut19_8), .EastIn(nOut20_7), .WestIn(nOut18_7), .ScanIn(nScanOut1224), .ScanOut(nScanOut1223), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_8), .NorthIn(nOut19_7), .SouthIn(nOut19_9), .EastIn(nOut20_8), .WestIn(nOut18_8), .ScanIn(nScanOut1225), .ScanOut(nScanOut1224), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_9), .NorthIn(nOut19_8), .SouthIn(nOut19_10), .EastIn(nOut20_9), .WestIn(nOut18_9), .ScanIn(nScanOut1226), .ScanOut(nScanOut1225), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_10), .NorthIn(nOut19_9), .SouthIn(nOut19_11), .EastIn(nOut20_10), .WestIn(nOut18_10), .ScanIn(nScanOut1227), .ScanOut(nScanOut1226), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_11), .NorthIn(nOut19_10), .SouthIn(nOut19_12), .EastIn(nOut20_11), .WestIn(nOut18_11), .ScanIn(nScanOut1228), .ScanOut(nScanOut1227), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_12), .NorthIn(nOut19_11), .SouthIn(nOut19_13), .EastIn(nOut20_12), .WestIn(nOut18_12), .ScanIn(nScanOut1229), .ScanOut(nScanOut1228), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_13), .NorthIn(nOut19_12), .SouthIn(nOut19_14), .EastIn(nOut20_13), .WestIn(nOut18_13), .ScanIn(nScanOut1230), .ScanOut(nScanOut1229), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_14), .NorthIn(nOut19_13), .SouthIn(nOut19_15), .EastIn(nOut20_14), .WestIn(nOut18_14), .ScanIn(nScanOut1231), .ScanOut(nScanOut1230), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_15), .NorthIn(nOut19_14), .SouthIn(nOut19_16), .EastIn(nOut20_15), .WestIn(nOut18_15), .ScanIn(nScanOut1232), .ScanOut(nScanOut1231), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_16), .NorthIn(nOut19_15), .SouthIn(nOut19_17), .EastIn(nOut20_16), .WestIn(nOut18_16), .ScanIn(nScanOut1233), .ScanOut(nScanOut1232), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_17), .NorthIn(nOut19_16), .SouthIn(nOut19_18), .EastIn(nOut20_17), .WestIn(nOut18_17), .ScanIn(nScanOut1234), .ScanOut(nScanOut1233), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_18), .NorthIn(nOut19_17), .SouthIn(nOut19_19), .EastIn(nOut20_18), .WestIn(nOut18_18), .ScanIn(nScanOut1235), .ScanOut(nScanOut1234), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_19), .NorthIn(nOut19_18), .SouthIn(nOut19_20), .EastIn(nOut20_19), .WestIn(nOut18_19), .ScanIn(nScanOut1236), .ScanOut(nScanOut1235), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_20), .NorthIn(nOut19_19), .SouthIn(nOut19_21), .EastIn(nOut20_20), .WestIn(nOut18_20), .ScanIn(nScanOut1237), .ScanOut(nScanOut1236), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_21), .NorthIn(nOut19_20), .SouthIn(nOut19_22), .EastIn(nOut20_21), .WestIn(nOut18_21), .ScanIn(nScanOut1238), .ScanOut(nScanOut1237), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_22), .NorthIn(nOut19_21), .SouthIn(nOut19_23), .EastIn(nOut20_22), .WestIn(nOut18_22), .ScanIn(nScanOut1239), .ScanOut(nScanOut1238), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_23), .NorthIn(nOut19_22), .SouthIn(nOut19_24), .EastIn(nOut20_23), .WestIn(nOut18_23), .ScanIn(nScanOut1240), .ScanOut(nScanOut1239), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_24), .NorthIn(nOut19_23), .SouthIn(nOut19_25), .EastIn(nOut20_24), .WestIn(nOut18_24), .ScanIn(nScanOut1241), .ScanOut(nScanOut1240), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_25), .NorthIn(nOut19_24), .SouthIn(nOut19_26), .EastIn(nOut20_25), .WestIn(nOut18_25), .ScanIn(nScanOut1242), .ScanOut(nScanOut1241), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_26), .NorthIn(nOut19_25), .SouthIn(nOut19_27), .EastIn(nOut20_26), .WestIn(nOut18_26), .ScanIn(nScanOut1243), .ScanOut(nScanOut1242), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_27), .NorthIn(nOut19_26), .SouthIn(nOut19_28), .EastIn(nOut20_27), .WestIn(nOut18_27), .ScanIn(nScanOut1244), .ScanOut(nScanOut1243), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_28), .NorthIn(nOut19_27), .SouthIn(nOut19_29), .EastIn(nOut20_28), .WestIn(nOut18_28), .ScanIn(nScanOut1245), .ScanOut(nScanOut1244), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_29), .NorthIn(nOut19_28), .SouthIn(nOut19_30), .EastIn(nOut20_29), .WestIn(nOut18_29), .ScanIn(nScanOut1246), .ScanOut(nScanOut1245), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_30), .NorthIn(nOut19_29), .SouthIn(nOut19_31), .EastIn(nOut20_30), .WestIn(nOut18_30), .ScanIn(nScanOut1247), .ScanOut(nScanOut1246), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_31), .NorthIn(nOut19_30), .SouthIn(nOut19_32), .EastIn(nOut20_31), .WestIn(nOut18_31), .ScanIn(nScanOut1248), .ScanOut(nScanOut1247), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_32), .NorthIn(nOut19_31), .SouthIn(nOut19_33), .EastIn(nOut20_32), .WestIn(nOut18_32), .ScanIn(nScanOut1249), .ScanOut(nScanOut1248), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_33), .NorthIn(nOut19_32), .SouthIn(nOut19_34), .EastIn(nOut20_33), .WestIn(nOut18_33), .ScanIn(nScanOut1250), .ScanOut(nScanOut1249), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_34), .NorthIn(nOut19_33), .SouthIn(nOut19_35), .EastIn(nOut20_34), .WestIn(nOut18_34), .ScanIn(nScanOut1251), .ScanOut(nScanOut1250), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_35), .NorthIn(nOut19_34), .SouthIn(nOut19_36), .EastIn(nOut20_35), .WestIn(nOut18_35), .ScanIn(nScanOut1252), .ScanOut(nScanOut1251), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_36), .NorthIn(nOut19_35), .SouthIn(nOut19_37), .EastIn(nOut20_36), .WestIn(nOut18_36), .ScanIn(nScanOut1253), .ScanOut(nScanOut1252), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_37), .NorthIn(nOut19_36), .SouthIn(nOut19_38), .EastIn(nOut20_37), .WestIn(nOut18_37), .ScanIn(nScanOut1254), .ScanOut(nScanOut1253), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_38), .NorthIn(nOut19_37), .SouthIn(nOut19_39), .EastIn(nOut20_38), .WestIn(nOut18_38), .ScanIn(nScanOut1255), .ScanOut(nScanOut1254), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_39), .NorthIn(nOut19_38), .SouthIn(nOut19_40), .EastIn(nOut20_39), .WestIn(nOut18_39), .ScanIn(nScanOut1256), .ScanOut(nScanOut1255), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1256 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_40), .NorthIn(nOut19_39), .SouthIn(nOut19_41), .EastIn(nOut20_40), .WestIn(nOut18_40), .ScanIn(nScanOut1257), .ScanOut(nScanOut1256), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1257 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_41), .NorthIn(nOut19_40), .SouthIn(nOut19_42), .EastIn(nOut20_41), .WestIn(nOut18_41), .ScanIn(nScanOut1258), .ScanOut(nScanOut1257), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1258 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_42), .NorthIn(nOut19_41), .SouthIn(nOut19_43), .EastIn(nOut20_42), .WestIn(nOut18_42), .ScanIn(nScanOut1259), .ScanOut(nScanOut1258), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1259 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_43), .NorthIn(nOut19_42), .SouthIn(nOut19_44), .EastIn(nOut20_43), .WestIn(nOut18_43), .ScanIn(nScanOut1260), .ScanOut(nScanOut1259), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1260 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_44), .NorthIn(nOut19_43), .SouthIn(nOut19_45), .EastIn(nOut20_44), .WestIn(nOut18_44), .ScanIn(nScanOut1261), .ScanOut(nScanOut1260), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1261 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_45), .NorthIn(nOut19_44), .SouthIn(nOut19_46), .EastIn(nOut20_45), .WestIn(nOut18_45), .ScanIn(nScanOut1262), .ScanOut(nScanOut1261), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1262 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_46), .NorthIn(nOut19_45), .SouthIn(nOut19_47), .EastIn(nOut20_46), .WestIn(nOut18_46), .ScanIn(nScanOut1263), .ScanOut(nScanOut1262), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1263 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_47), .NorthIn(nOut19_46), .SouthIn(nOut19_48), .EastIn(nOut20_47), .WestIn(nOut18_47), .ScanIn(nScanOut1264), .ScanOut(nScanOut1263), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1264 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_48), .NorthIn(nOut19_47), .SouthIn(nOut19_49), .EastIn(nOut20_48), .WestIn(nOut18_48), .ScanIn(nScanOut1265), .ScanOut(nScanOut1264), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1265 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_49), .NorthIn(nOut19_48), .SouthIn(nOut19_50), .EastIn(nOut20_49), .WestIn(nOut18_49), .ScanIn(nScanOut1266), .ScanOut(nScanOut1265), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1266 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_50), .NorthIn(nOut19_49), .SouthIn(nOut19_51), .EastIn(nOut20_50), .WestIn(nOut18_50), .ScanIn(nScanOut1267), .ScanOut(nScanOut1266), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1267 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_51), .NorthIn(nOut19_50), .SouthIn(nOut19_52), .EastIn(nOut20_51), .WestIn(nOut18_51), .ScanIn(nScanOut1268), .ScanOut(nScanOut1267), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1268 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_52), .NorthIn(nOut19_51), .SouthIn(nOut19_53), .EastIn(nOut20_52), .WestIn(nOut18_52), .ScanIn(nScanOut1269), .ScanOut(nScanOut1268), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1269 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_53), .NorthIn(nOut19_52), .SouthIn(nOut19_54), .EastIn(nOut20_53), .WestIn(nOut18_53), .ScanIn(nScanOut1270), .ScanOut(nScanOut1269), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1270 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_54), .NorthIn(nOut19_53), .SouthIn(nOut19_55), .EastIn(nOut20_54), .WestIn(nOut18_54), .ScanIn(nScanOut1271), .ScanOut(nScanOut1270), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1271 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_55), .NorthIn(nOut19_54), .SouthIn(nOut19_56), .EastIn(nOut20_55), .WestIn(nOut18_55), .ScanIn(nScanOut1272), .ScanOut(nScanOut1271), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1272 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_56), .NorthIn(nOut19_55), .SouthIn(nOut19_57), .EastIn(nOut20_56), .WestIn(nOut18_56), .ScanIn(nScanOut1273), .ScanOut(nScanOut1272), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1273 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_57), .NorthIn(nOut19_56), .SouthIn(nOut19_58), .EastIn(nOut20_57), .WestIn(nOut18_57), .ScanIn(nScanOut1274), .ScanOut(nScanOut1273), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1274 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_58), .NorthIn(nOut19_57), .SouthIn(nOut19_59), .EastIn(nOut20_58), .WestIn(nOut18_58), .ScanIn(nScanOut1275), .ScanOut(nScanOut1274), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1275 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_59), .NorthIn(nOut19_58), .SouthIn(nOut19_60), .EastIn(nOut20_59), .WestIn(nOut18_59), .ScanIn(nScanOut1276), .ScanOut(nScanOut1275), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1276 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_60), .NorthIn(nOut19_59), .SouthIn(nOut19_61), .EastIn(nOut20_60), .WestIn(nOut18_60), .ScanIn(nScanOut1277), .ScanOut(nScanOut1276), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1277 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_61), .NorthIn(nOut19_60), .SouthIn(nOut19_62), .EastIn(nOut20_61), .WestIn(nOut18_61), .ScanIn(nScanOut1278), .ScanOut(nScanOut1277), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1278 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut19_62), .NorthIn(nOut19_61), .SouthIn(nOut19_63), .EastIn(nOut20_62), .WestIn(nOut18_62), .ScanIn(nScanOut1279), .ScanOut(nScanOut1278), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1279 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut19_63), .ScanIn(nScanOut1280), .ScanOut(nScanOut1279), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1280 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut20_0), .ScanIn(nScanOut1281), .ScanOut(nScanOut1280), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1281 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_1), .NorthIn(nOut20_0), .SouthIn(nOut20_2), .EastIn(nOut21_1), .WestIn(nOut19_1), .ScanIn(nScanOut1282), .ScanOut(nScanOut1281), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1282 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_2), .NorthIn(nOut20_1), .SouthIn(nOut20_3), .EastIn(nOut21_2), .WestIn(nOut19_2), .ScanIn(nScanOut1283), .ScanOut(nScanOut1282), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1283 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_3), .NorthIn(nOut20_2), .SouthIn(nOut20_4), .EastIn(nOut21_3), .WestIn(nOut19_3), .ScanIn(nScanOut1284), .ScanOut(nScanOut1283), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1284 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_4), .NorthIn(nOut20_3), .SouthIn(nOut20_5), .EastIn(nOut21_4), .WestIn(nOut19_4), .ScanIn(nScanOut1285), .ScanOut(nScanOut1284), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1285 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_5), .NorthIn(nOut20_4), .SouthIn(nOut20_6), .EastIn(nOut21_5), .WestIn(nOut19_5), .ScanIn(nScanOut1286), .ScanOut(nScanOut1285), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1286 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_6), .NorthIn(nOut20_5), .SouthIn(nOut20_7), .EastIn(nOut21_6), .WestIn(nOut19_6), .ScanIn(nScanOut1287), .ScanOut(nScanOut1286), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1287 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_7), .NorthIn(nOut20_6), .SouthIn(nOut20_8), .EastIn(nOut21_7), .WestIn(nOut19_7), .ScanIn(nScanOut1288), .ScanOut(nScanOut1287), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1288 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_8), .NorthIn(nOut20_7), .SouthIn(nOut20_9), .EastIn(nOut21_8), .WestIn(nOut19_8), .ScanIn(nScanOut1289), .ScanOut(nScanOut1288), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1289 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_9), .NorthIn(nOut20_8), .SouthIn(nOut20_10), .EastIn(nOut21_9), .WestIn(nOut19_9), .ScanIn(nScanOut1290), .ScanOut(nScanOut1289), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1290 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_10), .NorthIn(nOut20_9), .SouthIn(nOut20_11), .EastIn(nOut21_10), .WestIn(nOut19_10), .ScanIn(nScanOut1291), .ScanOut(nScanOut1290), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1291 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_11), .NorthIn(nOut20_10), .SouthIn(nOut20_12), .EastIn(nOut21_11), .WestIn(nOut19_11), .ScanIn(nScanOut1292), .ScanOut(nScanOut1291), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1292 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_12), .NorthIn(nOut20_11), .SouthIn(nOut20_13), .EastIn(nOut21_12), .WestIn(nOut19_12), .ScanIn(nScanOut1293), .ScanOut(nScanOut1292), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1293 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_13), .NorthIn(nOut20_12), .SouthIn(nOut20_14), .EastIn(nOut21_13), .WestIn(nOut19_13), .ScanIn(nScanOut1294), .ScanOut(nScanOut1293), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1294 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_14), .NorthIn(nOut20_13), .SouthIn(nOut20_15), .EastIn(nOut21_14), .WestIn(nOut19_14), .ScanIn(nScanOut1295), .ScanOut(nScanOut1294), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1295 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_15), .NorthIn(nOut20_14), .SouthIn(nOut20_16), .EastIn(nOut21_15), .WestIn(nOut19_15), .ScanIn(nScanOut1296), .ScanOut(nScanOut1295), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1296 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_16), .NorthIn(nOut20_15), .SouthIn(nOut20_17), .EastIn(nOut21_16), .WestIn(nOut19_16), .ScanIn(nScanOut1297), .ScanOut(nScanOut1296), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1297 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_17), .NorthIn(nOut20_16), .SouthIn(nOut20_18), .EastIn(nOut21_17), .WestIn(nOut19_17), .ScanIn(nScanOut1298), .ScanOut(nScanOut1297), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1298 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_18), .NorthIn(nOut20_17), .SouthIn(nOut20_19), .EastIn(nOut21_18), .WestIn(nOut19_18), .ScanIn(nScanOut1299), .ScanOut(nScanOut1298), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1299 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_19), .NorthIn(nOut20_18), .SouthIn(nOut20_20), .EastIn(nOut21_19), .WestIn(nOut19_19), .ScanIn(nScanOut1300), .ScanOut(nScanOut1299), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1300 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_20), .NorthIn(nOut20_19), .SouthIn(nOut20_21), .EastIn(nOut21_20), .WestIn(nOut19_20), .ScanIn(nScanOut1301), .ScanOut(nScanOut1300), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1301 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_21), .NorthIn(nOut20_20), .SouthIn(nOut20_22), .EastIn(nOut21_21), .WestIn(nOut19_21), .ScanIn(nScanOut1302), .ScanOut(nScanOut1301), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1302 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_22), .NorthIn(nOut20_21), .SouthIn(nOut20_23), .EastIn(nOut21_22), .WestIn(nOut19_22), .ScanIn(nScanOut1303), .ScanOut(nScanOut1302), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1303 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_23), .NorthIn(nOut20_22), .SouthIn(nOut20_24), .EastIn(nOut21_23), .WestIn(nOut19_23), .ScanIn(nScanOut1304), .ScanOut(nScanOut1303), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1304 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_24), .NorthIn(nOut20_23), .SouthIn(nOut20_25), .EastIn(nOut21_24), .WestIn(nOut19_24), .ScanIn(nScanOut1305), .ScanOut(nScanOut1304), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1305 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_25), .NorthIn(nOut20_24), .SouthIn(nOut20_26), .EastIn(nOut21_25), .WestIn(nOut19_25), .ScanIn(nScanOut1306), .ScanOut(nScanOut1305), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1306 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_26), .NorthIn(nOut20_25), .SouthIn(nOut20_27), .EastIn(nOut21_26), .WestIn(nOut19_26), .ScanIn(nScanOut1307), .ScanOut(nScanOut1306), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1307 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_27), .NorthIn(nOut20_26), .SouthIn(nOut20_28), .EastIn(nOut21_27), .WestIn(nOut19_27), .ScanIn(nScanOut1308), .ScanOut(nScanOut1307), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1308 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_28), .NorthIn(nOut20_27), .SouthIn(nOut20_29), .EastIn(nOut21_28), .WestIn(nOut19_28), .ScanIn(nScanOut1309), .ScanOut(nScanOut1308), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1309 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_29), .NorthIn(nOut20_28), .SouthIn(nOut20_30), .EastIn(nOut21_29), .WestIn(nOut19_29), .ScanIn(nScanOut1310), .ScanOut(nScanOut1309), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1310 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_30), .NorthIn(nOut20_29), .SouthIn(nOut20_31), .EastIn(nOut21_30), .WestIn(nOut19_30), .ScanIn(nScanOut1311), .ScanOut(nScanOut1310), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1311 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_31), .NorthIn(nOut20_30), .SouthIn(nOut20_32), .EastIn(nOut21_31), .WestIn(nOut19_31), .ScanIn(nScanOut1312), .ScanOut(nScanOut1311), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1312 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_32), .NorthIn(nOut20_31), .SouthIn(nOut20_33), .EastIn(nOut21_32), .WestIn(nOut19_32), .ScanIn(nScanOut1313), .ScanOut(nScanOut1312), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1313 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_33), .NorthIn(nOut20_32), .SouthIn(nOut20_34), .EastIn(nOut21_33), .WestIn(nOut19_33), .ScanIn(nScanOut1314), .ScanOut(nScanOut1313), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1314 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_34), .NorthIn(nOut20_33), .SouthIn(nOut20_35), .EastIn(nOut21_34), .WestIn(nOut19_34), .ScanIn(nScanOut1315), .ScanOut(nScanOut1314), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1315 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_35), .NorthIn(nOut20_34), .SouthIn(nOut20_36), .EastIn(nOut21_35), .WestIn(nOut19_35), .ScanIn(nScanOut1316), .ScanOut(nScanOut1315), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1316 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_36), .NorthIn(nOut20_35), .SouthIn(nOut20_37), .EastIn(nOut21_36), .WestIn(nOut19_36), .ScanIn(nScanOut1317), .ScanOut(nScanOut1316), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1317 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_37), .NorthIn(nOut20_36), .SouthIn(nOut20_38), .EastIn(nOut21_37), .WestIn(nOut19_37), .ScanIn(nScanOut1318), .ScanOut(nScanOut1317), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1318 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_38), .NorthIn(nOut20_37), .SouthIn(nOut20_39), .EastIn(nOut21_38), .WestIn(nOut19_38), .ScanIn(nScanOut1319), .ScanOut(nScanOut1318), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1319 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_39), .NorthIn(nOut20_38), .SouthIn(nOut20_40), .EastIn(nOut21_39), .WestIn(nOut19_39), .ScanIn(nScanOut1320), .ScanOut(nScanOut1319), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1320 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_40), .NorthIn(nOut20_39), .SouthIn(nOut20_41), .EastIn(nOut21_40), .WestIn(nOut19_40), .ScanIn(nScanOut1321), .ScanOut(nScanOut1320), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1321 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_41), .NorthIn(nOut20_40), .SouthIn(nOut20_42), .EastIn(nOut21_41), .WestIn(nOut19_41), .ScanIn(nScanOut1322), .ScanOut(nScanOut1321), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1322 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_42), .NorthIn(nOut20_41), .SouthIn(nOut20_43), .EastIn(nOut21_42), .WestIn(nOut19_42), .ScanIn(nScanOut1323), .ScanOut(nScanOut1322), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1323 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_43), .NorthIn(nOut20_42), .SouthIn(nOut20_44), .EastIn(nOut21_43), .WestIn(nOut19_43), .ScanIn(nScanOut1324), .ScanOut(nScanOut1323), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1324 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_44), .NorthIn(nOut20_43), .SouthIn(nOut20_45), .EastIn(nOut21_44), .WestIn(nOut19_44), .ScanIn(nScanOut1325), .ScanOut(nScanOut1324), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1325 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_45), .NorthIn(nOut20_44), .SouthIn(nOut20_46), .EastIn(nOut21_45), .WestIn(nOut19_45), .ScanIn(nScanOut1326), .ScanOut(nScanOut1325), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1326 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_46), .NorthIn(nOut20_45), .SouthIn(nOut20_47), .EastIn(nOut21_46), .WestIn(nOut19_46), .ScanIn(nScanOut1327), .ScanOut(nScanOut1326), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1327 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_47), .NorthIn(nOut20_46), .SouthIn(nOut20_48), .EastIn(nOut21_47), .WestIn(nOut19_47), .ScanIn(nScanOut1328), .ScanOut(nScanOut1327), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1328 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_48), .NorthIn(nOut20_47), .SouthIn(nOut20_49), .EastIn(nOut21_48), .WestIn(nOut19_48), .ScanIn(nScanOut1329), .ScanOut(nScanOut1328), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1329 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_49), .NorthIn(nOut20_48), .SouthIn(nOut20_50), .EastIn(nOut21_49), .WestIn(nOut19_49), .ScanIn(nScanOut1330), .ScanOut(nScanOut1329), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1330 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_50), .NorthIn(nOut20_49), .SouthIn(nOut20_51), .EastIn(nOut21_50), .WestIn(nOut19_50), .ScanIn(nScanOut1331), .ScanOut(nScanOut1330), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1331 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_51), .NorthIn(nOut20_50), .SouthIn(nOut20_52), .EastIn(nOut21_51), .WestIn(nOut19_51), .ScanIn(nScanOut1332), .ScanOut(nScanOut1331), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1332 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_52), .NorthIn(nOut20_51), .SouthIn(nOut20_53), .EastIn(nOut21_52), .WestIn(nOut19_52), .ScanIn(nScanOut1333), .ScanOut(nScanOut1332), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1333 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_53), .NorthIn(nOut20_52), .SouthIn(nOut20_54), .EastIn(nOut21_53), .WestIn(nOut19_53), .ScanIn(nScanOut1334), .ScanOut(nScanOut1333), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1334 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_54), .NorthIn(nOut20_53), .SouthIn(nOut20_55), .EastIn(nOut21_54), .WestIn(nOut19_54), .ScanIn(nScanOut1335), .ScanOut(nScanOut1334), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1335 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_55), .NorthIn(nOut20_54), .SouthIn(nOut20_56), .EastIn(nOut21_55), .WestIn(nOut19_55), .ScanIn(nScanOut1336), .ScanOut(nScanOut1335), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1336 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_56), .NorthIn(nOut20_55), .SouthIn(nOut20_57), .EastIn(nOut21_56), .WestIn(nOut19_56), .ScanIn(nScanOut1337), .ScanOut(nScanOut1336), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1337 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_57), .NorthIn(nOut20_56), .SouthIn(nOut20_58), .EastIn(nOut21_57), .WestIn(nOut19_57), .ScanIn(nScanOut1338), .ScanOut(nScanOut1337), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1338 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_58), .NorthIn(nOut20_57), .SouthIn(nOut20_59), .EastIn(nOut21_58), .WestIn(nOut19_58), .ScanIn(nScanOut1339), .ScanOut(nScanOut1338), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1339 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_59), .NorthIn(nOut20_58), .SouthIn(nOut20_60), .EastIn(nOut21_59), .WestIn(nOut19_59), .ScanIn(nScanOut1340), .ScanOut(nScanOut1339), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1340 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_60), .NorthIn(nOut20_59), .SouthIn(nOut20_61), .EastIn(nOut21_60), .WestIn(nOut19_60), .ScanIn(nScanOut1341), .ScanOut(nScanOut1340), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1341 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_61), .NorthIn(nOut20_60), .SouthIn(nOut20_62), .EastIn(nOut21_61), .WestIn(nOut19_61), .ScanIn(nScanOut1342), .ScanOut(nScanOut1341), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1342 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut20_62), .NorthIn(nOut20_61), .SouthIn(nOut20_63), .EastIn(nOut21_62), .WestIn(nOut19_62), .ScanIn(nScanOut1343), .ScanOut(nScanOut1342), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1343 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut20_63), .ScanIn(nScanOut1344), .ScanOut(nScanOut1343), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1344 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut21_0), .ScanIn(nScanOut1345), .ScanOut(nScanOut1344), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1345 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_1), .NorthIn(nOut21_0), .SouthIn(nOut21_2), .EastIn(nOut22_1), .WestIn(nOut20_1), .ScanIn(nScanOut1346), .ScanOut(nScanOut1345), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1346 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_2), .NorthIn(nOut21_1), .SouthIn(nOut21_3), .EastIn(nOut22_2), .WestIn(nOut20_2), .ScanIn(nScanOut1347), .ScanOut(nScanOut1346), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1347 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_3), .NorthIn(nOut21_2), .SouthIn(nOut21_4), .EastIn(nOut22_3), .WestIn(nOut20_3), .ScanIn(nScanOut1348), .ScanOut(nScanOut1347), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1348 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_4), .NorthIn(nOut21_3), .SouthIn(nOut21_5), .EastIn(nOut22_4), .WestIn(nOut20_4), .ScanIn(nScanOut1349), .ScanOut(nScanOut1348), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1349 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_5), .NorthIn(nOut21_4), .SouthIn(nOut21_6), .EastIn(nOut22_5), .WestIn(nOut20_5), .ScanIn(nScanOut1350), .ScanOut(nScanOut1349), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1350 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_6), .NorthIn(nOut21_5), .SouthIn(nOut21_7), .EastIn(nOut22_6), .WestIn(nOut20_6), .ScanIn(nScanOut1351), .ScanOut(nScanOut1350), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1351 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_7), .NorthIn(nOut21_6), .SouthIn(nOut21_8), .EastIn(nOut22_7), .WestIn(nOut20_7), .ScanIn(nScanOut1352), .ScanOut(nScanOut1351), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1352 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_8), .NorthIn(nOut21_7), .SouthIn(nOut21_9), .EastIn(nOut22_8), .WestIn(nOut20_8), .ScanIn(nScanOut1353), .ScanOut(nScanOut1352), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1353 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_9), .NorthIn(nOut21_8), .SouthIn(nOut21_10), .EastIn(nOut22_9), .WestIn(nOut20_9), .ScanIn(nScanOut1354), .ScanOut(nScanOut1353), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1354 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_10), .NorthIn(nOut21_9), .SouthIn(nOut21_11), .EastIn(nOut22_10), .WestIn(nOut20_10), .ScanIn(nScanOut1355), .ScanOut(nScanOut1354), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1355 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_11), .NorthIn(nOut21_10), .SouthIn(nOut21_12), .EastIn(nOut22_11), .WestIn(nOut20_11), .ScanIn(nScanOut1356), .ScanOut(nScanOut1355), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1356 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_12), .NorthIn(nOut21_11), .SouthIn(nOut21_13), .EastIn(nOut22_12), .WestIn(nOut20_12), .ScanIn(nScanOut1357), .ScanOut(nScanOut1356), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1357 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_13), .NorthIn(nOut21_12), .SouthIn(nOut21_14), .EastIn(nOut22_13), .WestIn(nOut20_13), .ScanIn(nScanOut1358), .ScanOut(nScanOut1357), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1358 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_14), .NorthIn(nOut21_13), .SouthIn(nOut21_15), .EastIn(nOut22_14), .WestIn(nOut20_14), .ScanIn(nScanOut1359), .ScanOut(nScanOut1358), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1359 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_15), .NorthIn(nOut21_14), .SouthIn(nOut21_16), .EastIn(nOut22_15), .WestIn(nOut20_15), .ScanIn(nScanOut1360), .ScanOut(nScanOut1359), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1360 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_16), .NorthIn(nOut21_15), .SouthIn(nOut21_17), .EastIn(nOut22_16), .WestIn(nOut20_16), .ScanIn(nScanOut1361), .ScanOut(nScanOut1360), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1361 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_17), .NorthIn(nOut21_16), .SouthIn(nOut21_18), .EastIn(nOut22_17), .WestIn(nOut20_17), .ScanIn(nScanOut1362), .ScanOut(nScanOut1361), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1362 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_18), .NorthIn(nOut21_17), .SouthIn(nOut21_19), .EastIn(nOut22_18), .WestIn(nOut20_18), .ScanIn(nScanOut1363), .ScanOut(nScanOut1362), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1363 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_19), .NorthIn(nOut21_18), .SouthIn(nOut21_20), .EastIn(nOut22_19), .WestIn(nOut20_19), .ScanIn(nScanOut1364), .ScanOut(nScanOut1363), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1364 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_20), .NorthIn(nOut21_19), .SouthIn(nOut21_21), .EastIn(nOut22_20), .WestIn(nOut20_20), .ScanIn(nScanOut1365), .ScanOut(nScanOut1364), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1365 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_21), .NorthIn(nOut21_20), .SouthIn(nOut21_22), .EastIn(nOut22_21), .WestIn(nOut20_21), .ScanIn(nScanOut1366), .ScanOut(nScanOut1365), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1366 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_22), .NorthIn(nOut21_21), .SouthIn(nOut21_23), .EastIn(nOut22_22), .WestIn(nOut20_22), .ScanIn(nScanOut1367), .ScanOut(nScanOut1366), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1367 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_23), .NorthIn(nOut21_22), .SouthIn(nOut21_24), .EastIn(nOut22_23), .WestIn(nOut20_23), .ScanIn(nScanOut1368), .ScanOut(nScanOut1367), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1368 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_24), .NorthIn(nOut21_23), .SouthIn(nOut21_25), .EastIn(nOut22_24), .WestIn(nOut20_24), .ScanIn(nScanOut1369), .ScanOut(nScanOut1368), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1369 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_25), .NorthIn(nOut21_24), .SouthIn(nOut21_26), .EastIn(nOut22_25), .WestIn(nOut20_25), .ScanIn(nScanOut1370), .ScanOut(nScanOut1369), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1370 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_26), .NorthIn(nOut21_25), .SouthIn(nOut21_27), .EastIn(nOut22_26), .WestIn(nOut20_26), .ScanIn(nScanOut1371), .ScanOut(nScanOut1370), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1371 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_27), .NorthIn(nOut21_26), .SouthIn(nOut21_28), .EastIn(nOut22_27), .WestIn(nOut20_27), .ScanIn(nScanOut1372), .ScanOut(nScanOut1371), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1372 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_28), .NorthIn(nOut21_27), .SouthIn(nOut21_29), .EastIn(nOut22_28), .WestIn(nOut20_28), .ScanIn(nScanOut1373), .ScanOut(nScanOut1372), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1373 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_29), .NorthIn(nOut21_28), .SouthIn(nOut21_30), .EastIn(nOut22_29), .WestIn(nOut20_29), .ScanIn(nScanOut1374), .ScanOut(nScanOut1373), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1374 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_30), .NorthIn(nOut21_29), .SouthIn(nOut21_31), .EastIn(nOut22_30), .WestIn(nOut20_30), .ScanIn(nScanOut1375), .ScanOut(nScanOut1374), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1375 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_31), .NorthIn(nOut21_30), .SouthIn(nOut21_32), .EastIn(nOut22_31), .WestIn(nOut20_31), .ScanIn(nScanOut1376), .ScanOut(nScanOut1375), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1376 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_32), .NorthIn(nOut21_31), .SouthIn(nOut21_33), .EastIn(nOut22_32), .WestIn(nOut20_32), .ScanIn(nScanOut1377), .ScanOut(nScanOut1376), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1377 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_33), .NorthIn(nOut21_32), .SouthIn(nOut21_34), .EastIn(nOut22_33), .WestIn(nOut20_33), .ScanIn(nScanOut1378), .ScanOut(nScanOut1377), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1378 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_34), .NorthIn(nOut21_33), .SouthIn(nOut21_35), .EastIn(nOut22_34), .WestIn(nOut20_34), .ScanIn(nScanOut1379), .ScanOut(nScanOut1378), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1379 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_35), .NorthIn(nOut21_34), .SouthIn(nOut21_36), .EastIn(nOut22_35), .WestIn(nOut20_35), .ScanIn(nScanOut1380), .ScanOut(nScanOut1379), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1380 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_36), .NorthIn(nOut21_35), .SouthIn(nOut21_37), .EastIn(nOut22_36), .WestIn(nOut20_36), .ScanIn(nScanOut1381), .ScanOut(nScanOut1380), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1381 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_37), .NorthIn(nOut21_36), .SouthIn(nOut21_38), .EastIn(nOut22_37), .WestIn(nOut20_37), .ScanIn(nScanOut1382), .ScanOut(nScanOut1381), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1382 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_38), .NorthIn(nOut21_37), .SouthIn(nOut21_39), .EastIn(nOut22_38), .WestIn(nOut20_38), .ScanIn(nScanOut1383), .ScanOut(nScanOut1382), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1383 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_39), .NorthIn(nOut21_38), .SouthIn(nOut21_40), .EastIn(nOut22_39), .WestIn(nOut20_39), .ScanIn(nScanOut1384), .ScanOut(nScanOut1383), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1384 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_40), .NorthIn(nOut21_39), .SouthIn(nOut21_41), .EastIn(nOut22_40), .WestIn(nOut20_40), .ScanIn(nScanOut1385), .ScanOut(nScanOut1384), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1385 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_41), .NorthIn(nOut21_40), .SouthIn(nOut21_42), .EastIn(nOut22_41), .WestIn(nOut20_41), .ScanIn(nScanOut1386), .ScanOut(nScanOut1385), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1386 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_42), .NorthIn(nOut21_41), .SouthIn(nOut21_43), .EastIn(nOut22_42), .WestIn(nOut20_42), .ScanIn(nScanOut1387), .ScanOut(nScanOut1386), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1387 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_43), .NorthIn(nOut21_42), .SouthIn(nOut21_44), .EastIn(nOut22_43), .WestIn(nOut20_43), .ScanIn(nScanOut1388), .ScanOut(nScanOut1387), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1388 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_44), .NorthIn(nOut21_43), .SouthIn(nOut21_45), .EastIn(nOut22_44), .WestIn(nOut20_44), .ScanIn(nScanOut1389), .ScanOut(nScanOut1388), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1389 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_45), .NorthIn(nOut21_44), .SouthIn(nOut21_46), .EastIn(nOut22_45), .WestIn(nOut20_45), .ScanIn(nScanOut1390), .ScanOut(nScanOut1389), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1390 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_46), .NorthIn(nOut21_45), .SouthIn(nOut21_47), .EastIn(nOut22_46), .WestIn(nOut20_46), .ScanIn(nScanOut1391), .ScanOut(nScanOut1390), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1391 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_47), .NorthIn(nOut21_46), .SouthIn(nOut21_48), .EastIn(nOut22_47), .WestIn(nOut20_47), .ScanIn(nScanOut1392), .ScanOut(nScanOut1391), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1392 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_48), .NorthIn(nOut21_47), .SouthIn(nOut21_49), .EastIn(nOut22_48), .WestIn(nOut20_48), .ScanIn(nScanOut1393), .ScanOut(nScanOut1392), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1393 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_49), .NorthIn(nOut21_48), .SouthIn(nOut21_50), .EastIn(nOut22_49), .WestIn(nOut20_49), .ScanIn(nScanOut1394), .ScanOut(nScanOut1393), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1394 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_50), .NorthIn(nOut21_49), .SouthIn(nOut21_51), .EastIn(nOut22_50), .WestIn(nOut20_50), .ScanIn(nScanOut1395), .ScanOut(nScanOut1394), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1395 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_51), .NorthIn(nOut21_50), .SouthIn(nOut21_52), .EastIn(nOut22_51), .WestIn(nOut20_51), .ScanIn(nScanOut1396), .ScanOut(nScanOut1395), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1396 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_52), .NorthIn(nOut21_51), .SouthIn(nOut21_53), .EastIn(nOut22_52), .WestIn(nOut20_52), .ScanIn(nScanOut1397), .ScanOut(nScanOut1396), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1397 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_53), .NorthIn(nOut21_52), .SouthIn(nOut21_54), .EastIn(nOut22_53), .WestIn(nOut20_53), .ScanIn(nScanOut1398), .ScanOut(nScanOut1397), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1398 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_54), .NorthIn(nOut21_53), .SouthIn(nOut21_55), .EastIn(nOut22_54), .WestIn(nOut20_54), .ScanIn(nScanOut1399), .ScanOut(nScanOut1398), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1399 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_55), .NorthIn(nOut21_54), .SouthIn(nOut21_56), .EastIn(nOut22_55), .WestIn(nOut20_55), .ScanIn(nScanOut1400), .ScanOut(nScanOut1399), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1400 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_56), .NorthIn(nOut21_55), .SouthIn(nOut21_57), .EastIn(nOut22_56), .WestIn(nOut20_56), .ScanIn(nScanOut1401), .ScanOut(nScanOut1400), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1401 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_57), .NorthIn(nOut21_56), .SouthIn(nOut21_58), .EastIn(nOut22_57), .WestIn(nOut20_57), .ScanIn(nScanOut1402), .ScanOut(nScanOut1401), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1402 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_58), .NorthIn(nOut21_57), .SouthIn(nOut21_59), .EastIn(nOut22_58), .WestIn(nOut20_58), .ScanIn(nScanOut1403), .ScanOut(nScanOut1402), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1403 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_59), .NorthIn(nOut21_58), .SouthIn(nOut21_60), .EastIn(nOut22_59), .WestIn(nOut20_59), .ScanIn(nScanOut1404), .ScanOut(nScanOut1403), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1404 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_60), .NorthIn(nOut21_59), .SouthIn(nOut21_61), .EastIn(nOut22_60), .WestIn(nOut20_60), .ScanIn(nScanOut1405), .ScanOut(nScanOut1404), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1405 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_61), .NorthIn(nOut21_60), .SouthIn(nOut21_62), .EastIn(nOut22_61), .WestIn(nOut20_61), .ScanIn(nScanOut1406), .ScanOut(nScanOut1405), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1406 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut21_62), .NorthIn(nOut21_61), .SouthIn(nOut21_63), .EastIn(nOut22_62), .WestIn(nOut20_62), .ScanIn(nScanOut1407), .ScanOut(nScanOut1406), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1407 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut21_63), .ScanIn(nScanOut1408), .ScanOut(nScanOut1407), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1408 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut22_0), .ScanIn(nScanOut1409), .ScanOut(nScanOut1408), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1409 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_1), .NorthIn(nOut22_0), .SouthIn(nOut22_2), .EastIn(nOut23_1), .WestIn(nOut21_1), .ScanIn(nScanOut1410), .ScanOut(nScanOut1409), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1410 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_2), .NorthIn(nOut22_1), .SouthIn(nOut22_3), .EastIn(nOut23_2), .WestIn(nOut21_2), .ScanIn(nScanOut1411), .ScanOut(nScanOut1410), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1411 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_3), .NorthIn(nOut22_2), .SouthIn(nOut22_4), .EastIn(nOut23_3), .WestIn(nOut21_3), .ScanIn(nScanOut1412), .ScanOut(nScanOut1411), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1412 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_4), .NorthIn(nOut22_3), .SouthIn(nOut22_5), .EastIn(nOut23_4), .WestIn(nOut21_4), .ScanIn(nScanOut1413), .ScanOut(nScanOut1412), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1413 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_5), .NorthIn(nOut22_4), .SouthIn(nOut22_6), .EastIn(nOut23_5), .WestIn(nOut21_5), .ScanIn(nScanOut1414), .ScanOut(nScanOut1413), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1414 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_6), .NorthIn(nOut22_5), .SouthIn(nOut22_7), .EastIn(nOut23_6), .WestIn(nOut21_6), .ScanIn(nScanOut1415), .ScanOut(nScanOut1414), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1415 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_7), .NorthIn(nOut22_6), .SouthIn(nOut22_8), .EastIn(nOut23_7), .WestIn(nOut21_7), .ScanIn(nScanOut1416), .ScanOut(nScanOut1415), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1416 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_8), .NorthIn(nOut22_7), .SouthIn(nOut22_9), .EastIn(nOut23_8), .WestIn(nOut21_8), .ScanIn(nScanOut1417), .ScanOut(nScanOut1416), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1417 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_9), .NorthIn(nOut22_8), .SouthIn(nOut22_10), .EastIn(nOut23_9), .WestIn(nOut21_9), .ScanIn(nScanOut1418), .ScanOut(nScanOut1417), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1418 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_10), .NorthIn(nOut22_9), .SouthIn(nOut22_11), .EastIn(nOut23_10), .WestIn(nOut21_10), .ScanIn(nScanOut1419), .ScanOut(nScanOut1418), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1419 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_11), .NorthIn(nOut22_10), .SouthIn(nOut22_12), .EastIn(nOut23_11), .WestIn(nOut21_11), .ScanIn(nScanOut1420), .ScanOut(nScanOut1419), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1420 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_12), .NorthIn(nOut22_11), .SouthIn(nOut22_13), .EastIn(nOut23_12), .WestIn(nOut21_12), .ScanIn(nScanOut1421), .ScanOut(nScanOut1420), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1421 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_13), .NorthIn(nOut22_12), .SouthIn(nOut22_14), .EastIn(nOut23_13), .WestIn(nOut21_13), .ScanIn(nScanOut1422), .ScanOut(nScanOut1421), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1422 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_14), .NorthIn(nOut22_13), .SouthIn(nOut22_15), .EastIn(nOut23_14), .WestIn(nOut21_14), .ScanIn(nScanOut1423), .ScanOut(nScanOut1422), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1423 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_15), .NorthIn(nOut22_14), .SouthIn(nOut22_16), .EastIn(nOut23_15), .WestIn(nOut21_15), .ScanIn(nScanOut1424), .ScanOut(nScanOut1423), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1424 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_16), .NorthIn(nOut22_15), .SouthIn(nOut22_17), .EastIn(nOut23_16), .WestIn(nOut21_16), .ScanIn(nScanOut1425), .ScanOut(nScanOut1424), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1425 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_17), .NorthIn(nOut22_16), .SouthIn(nOut22_18), .EastIn(nOut23_17), .WestIn(nOut21_17), .ScanIn(nScanOut1426), .ScanOut(nScanOut1425), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1426 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_18), .NorthIn(nOut22_17), .SouthIn(nOut22_19), .EastIn(nOut23_18), .WestIn(nOut21_18), .ScanIn(nScanOut1427), .ScanOut(nScanOut1426), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1427 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_19), .NorthIn(nOut22_18), .SouthIn(nOut22_20), .EastIn(nOut23_19), .WestIn(nOut21_19), .ScanIn(nScanOut1428), .ScanOut(nScanOut1427), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1428 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_20), .NorthIn(nOut22_19), .SouthIn(nOut22_21), .EastIn(nOut23_20), .WestIn(nOut21_20), .ScanIn(nScanOut1429), .ScanOut(nScanOut1428), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1429 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_21), .NorthIn(nOut22_20), .SouthIn(nOut22_22), .EastIn(nOut23_21), .WestIn(nOut21_21), .ScanIn(nScanOut1430), .ScanOut(nScanOut1429), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1430 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_22), .NorthIn(nOut22_21), .SouthIn(nOut22_23), .EastIn(nOut23_22), .WestIn(nOut21_22), .ScanIn(nScanOut1431), .ScanOut(nScanOut1430), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1431 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_23), .NorthIn(nOut22_22), .SouthIn(nOut22_24), .EastIn(nOut23_23), .WestIn(nOut21_23), .ScanIn(nScanOut1432), .ScanOut(nScanOut1431), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1432 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_24), .NorthIn(nOut22_23), .SouthIn(nOut22_25), .EastIn(nOut23_24), .WestIn(nOut21_24), .ScanIn(nScanOut1433), .ScanOut(nScanOut1432), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1433 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_25), .NorthIn(nOut22_24), .SouthIn(nOut22_26), .EastIn(nOut23_25), .WestIn(nOut21_25), .ScanIn(nScanOut1434), .ScanOut(nScanOut1433), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1434 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_26), .NorthIn(nOut22_25), .SouthIn(nOut22_27), .EastIn(nOut23_26), .WestIn(nOut21_26), .ScanIn(nScanOut1435), .ScanOut(nScanOut1434), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1435 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_27), .NorthIn(nOut22_26), .SouthIn(nOut22_28), .EastIn(nOut23_27), .WestIn(nOut21_27), .ScanIn(nScanOut1436), .ScanOut(nScanOut1435), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1436 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_28), .NorthIn(nOut22_27), .SouthIn(nOut22_29), .EastIn(nOut23_28), .WestIn(nOut21_28), .ScanIn(nScanOut1437), .ScanOut(nScanOut1436), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1437 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_29), .NorthIn(nOut22_28), .SouthIn(nOut22_30), .EastIn(nOut23_29), .WestIn(nOut21_29), .ScanIn(nScanOut1438), .ScanOut(nScanOut1437), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1438 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_30), .NorthIn(nOut22_29), .SouthIn(nOut22_31), .EastIn(nOut23_30), .WestIn(nOut21_30), .ScanIn(nScanOut1439), .ScanOut(nScanOut1438), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1439 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_31), .NorthIn(nOut22_30), .SouthIn(nOut22_32), .EastIn(nOut23_31), .WestIn(nOut21_31), .ScanIn(nScanOut1440), .ScanOut(nScanOut1439), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1440 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_32), .NorthIn(nOut22_31), .SouthIn(nOut22_33), .EastIn(nOut23_32), .WestIn(nOut21_32), .ScanIn(nScanOut1441), .ScanOut(nScanOut1440), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1441 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_33), .NorthIn(nOut22_32), .SouthIn(nOut22_34), .EastIn(nOut23_33), .WestIn(nOut21_33), .ScanIn(nScanOut1442), .ScanOut(nScanOut1441), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1442 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_34), .NorthIn(nOut22_33), .SouthIn(nOut22_35), .EastIn(nOut23_34), .WestIn(nOut21_34), .ScanIn(nScanOut1443), .ScanOut(nScanOut1442), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1443 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_35), .NorthIn(nOut22_34), .SouthIn(nOut22_36), .EastIn(nOut23_35), .WestIn(nOut21_35), .ScanIn(nScanOut1444), .ScanOut(nScanOut1443), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1444 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_36), .NorthIn(nOut22_35), .SouthIn(nOut22_37), .EastIn(nOut23_36), .WestIn(nOut21_36), .ScanIn(nScanOut1445), .ScanOut(nScanOut1444), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1445 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_37), .NorthIn(nOut22_36), .SouthIn(nOut22_38), .EastIn(nOut23_37), .WestIn(nOut21_37), .ScanIn(nScanOut1446), .ScanOut(nScanOut1445), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1446 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_38), .NorthIn(nOut22_37), .SouthIn(nOut22_39), .EastIn(nOut23_38), .WestIn(nOut21_38), .ScanIn(nScanOut1447), .ScanOut(nScanOut1446), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1447 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_39), .NorthIn(nOut22_38), .SouthIn(nOut22_40), .EastIn(nOut23_39), .WestIn(nOut21_39), .ScanIn(nScanOut1448), .ScanOut(nScanOut1447), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1448 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_40), .NorthIn(nOut22_39), .SouthIn(nOut22_41), .EastIn(nOut23_40), .WestIn(nOut21_40), .ScanIn(nScanOut1449), .ScanOut(nScanOut1448), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1449 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_41), .NorthIn(nOut22_40), .SouthIn(nOut22_42), .EastIn(nOut23_41), .WestIn(nOut21_41), .ScanIn(nScanOut1450), .ScanOut(nScanOut1449), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1450 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_42), .NorthIn(nOut22_41), .SouthIn(nOut22_43), .EastIn(nOut23_42), .WestIn(nOut21_42), .ScanIn(nScanOut1451), .ScanOut(nScanOut1450), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1451 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_43), .NorthIn(nOut22_42), .SouthIn(nOut22_44), .EastIn(nOut23_43), .WestIn(nOut21_43), .ScanIn(nScanOut1452), .ScanOut(nScanOut1451), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1452 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_44), .NorthIn(nOut22_43), .SouthIn(nOut22_45), .EastIn(nOut23_44), .WestIn(nOut21_44), .ScanIn(nScanOut1453), .ScanOut(nScanOut1452), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1453 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_45), .NorthIn(nOut22_44), .SouthIn(nOut22_46), .EastIn(nOut23_45), .WestIn(nOut21_45), .ScanIn(nScanOut1454), .ScanOut(nScanOut1453), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1454 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_46), .NorthIn(nOut22_45), .SouthIn(nOut22_47), .EastIn(nOut23_46), .WestIn(nOut21_46), .ScanIn(nScanOut1455), .ScanOut(nScanOut1454), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1455 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_47), .NorthIn(nOut22_46), .SouthIn(nOut22_48), .EastIn(nOut23_47), .WestIn(nOut21_47), .ScanIn(nScanOut1456), .ScanOut(nScanOut1455), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1456 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_48), .NorthIn(nOut22_47), .SouthIn(nOut22_49), .EastIn(nOut23_48), .WestIn(nOut21_48), .ScanIn(nScanOut1457), .ScanOut(nScanOut1456), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1457 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_49), .NorthIn(nOut22_48), .SouthIn(nOut22_50), .EastIn(nOut23_49), .WestIn(nOut21_49), .ScanIn(nScanOut1458), .ScanOut(nScanOut1457), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1458 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_50), .NorthIn(nOut22_49), .SouthIn(nOut22_51), .EastIn(nOut23_50), .WestIn(nOut21_50), .ScanIn(nScanOut1459), .ScanOut(nScanOut1458), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1459 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_51), .NorthIn(nOut22_50), .SouthIn(nOut22_52), .EastIn(nOut23_51), .WestIn(nOut21_51), .ScanIn(nScanOut1460), .ScanOut(nScanOut1459), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1460 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_52), .NorthIn(nOut22_51), .SouthIn(nOut22_53), .EastIn(nOut23_52), .WestIn(nOut21_52), .ScanIn(nScanOut1461), .ScanOut(nScanOut1460), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1461 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_53), .NorthIn(nOut22_52), .SouthIn(nOut22_54), .EastIn(nOut23_53), .WestIn(nOut21_53), .ScanIn(nScanOut1462), .ScanOut(nScanOut1461), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1462 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_54), .NorthIn(nOut22_53), .SouthIn(nOut22_55), .EastIn(nOut23_54), .WestIn(nOut21_54), .ScanIn(nScanOut1463), .ScanOut(nScanOut1462), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1463 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_55), .NorthIn(nOut22_54), .SouthIn(nOut22_56), .EastIn(nOut23_55), .WestIn(nOut21_55), .ScanIn(nScanOut1464), .ScanOut(nScanOut1463), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1464 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_56), .NorthIn(nOut22_55), .SouthIn(nOut22_57), .EastIn(nOut23_56), .WestIn(nOut21_56), .ScanIn(nScanOut1465), .ScanOut(nScanOut1464), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1465 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_57), .NorthIn(nOut22_56), .SouthIn(nOut22_58), .EastIn(nOut23_57), .WestIn(nOut21_57), .ScanIn(nScanOut1466), .ScanOut(nScanOut1465), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1466 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_58), .NorthIn(nOut22_57), .SouthIn(nOut22_59), .EastIn(nOut23_58), .WestIn(nOut21_58), .ScanIn(nScanOut1467), .ScanOut(nScanOut1466), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1467 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_59), .NorthIn(nOut22_58), .SouthIn(nOut22_60), .EastIn(nOut23_59), .WestIn(nOut21_59), .ScanIn(nScanOut1468), .ScanOut(nScanOut1467), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1468 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_60), .NorthIn(nOut22_59), .SouthIn(nOut22_61), .EastIn(nOut23_60), .WestIn(nOut21_60), .ScanIn(nScanOut1469), .ScanOut(nScanOut1468), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1469 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_61), .NorthIn(nOut22_60), .SouthIn(nOut22_62), .EastIn(nOut23_61), .WestIn(nOut21_61), .ScanIn(nScanOut1470), .ScanOut(nScanOut1469), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1470 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut22_62), .NorthIn(nOut22_61), .SouthIn(nOut22_63), .EastIn(nOut23_62), .WestIn(nOut21_62), .ScanIn(nScanOut1471), .ScanOut(nScanOut1470), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1471 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut22_63), .ScanIn(nScanOut1472), .ScanOut(nScanOut1471), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1472 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut23_0), .ScanIn(nScanOut1473), .ScanOut(nScanOut1472), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1473 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_1), .NorthIn(nOut23_0), .SouthIn(nOut23_2), .EastIn(nOut24_1), .WestIn(nOut22_1), .ScanIn(nScanOut1474), .ScanOut(nScanOut1473), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1474 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_2), .NorthIn(nOut23_1), .SouthIn(nOut23_3), .EastIn(nOut24_2), .WestIn(nOut22_2), .ScanIn(nScanOut1475), .ScanOut(nScanOut1474), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1475 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_3), .NorthIn(nOut23_2), .SouthIn(nOut23_4), .EastIn(nOut24_3), .WestIn(nOut22_3), .ScanIn(nScanOut1476), .ScanOut(nScanOut1475), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1476 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_4), .NorthIn(nOut23_3), .SouthIn(nOut23_5), .EastIn(nOut24_4), .WestIn(nOut22_4), .ScanIn(nScanOut1477), .ScanOut(nScanOut1476), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1477 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_5), .NorthIn(nOut23_4), .SouthIn(nOut23_6), .EastIn(nOut24_5), .WestIn(nOut22_5), .ScanIn(nScanOut1478), .ScanOut(nScanOut1477), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1478 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_6), .NorthIn(nOut23_5), .SouthIn(nOut23_7), .EastIn(nOut24_6), .WestIn(nOut22_6), .ScanIn(nScanOut1479), .ScanOut(nScanOut1478), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1479 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_7), .NorthIn(nOut23_6), .SouthIn(nOut23_8), .EastIn(nOut24_7), .WestIn(nOut22_7), .ScanIn(nScanOut1480), .ScanOut(nScanOut1479), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1480 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_8), .NorthIn(nOut23_7), .SouthIn(nOut23_9), .EastIn(nOut24_8), .WestIn(nOut22_8), .ScanIn(nScanOut1481), .ScanOut(nScanOut1480), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1481 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_9), .NorthIn(nOut23_8), .SouthIn(nOut23_10), .EastIn(nOut24_9), .WestIn(nOut22_9), .ScanIn(nScanOut1482), .ScanOut(nScanOut1481), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1482 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_10), .NorthIn(nOut23_9), .SouthIn(nOut23_11), .EastIn(nOut24_10), .WestIn(nOut22_10), .ScanIn(nScanOut1483), .ScanOut(nScanOut1482), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1483 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_11), .NorthIn(nOut23_10), .SouthIn(nOut23_12), .EastIn(nOut24_11), .WestIn(nOut22_11), .ScanIn(nScanOut1484), .ScanOut(nScanOut1483), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1484 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_12), .NorthIn(nOut23_11), .SouthIn(nOut23_13), .EastIn(nOut24_12), .WestIn(nOut22_12), .ScanIn(nScanOut1485), .ScanOut(nScanOut1484), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1485 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_13), .NorthIn(nOut23_12), .SouthIn(nOut23_14), .EastIn(nOut24_13), .WestIn(nOut22_13), .ScanIn(nScanOut1486), .ScanOut(nScanOut1485), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1486 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_14), .NorthIn(nOut23_13), .SouthIn(nOut23_15), .EastIn(nOut24_14), .WestIn(nOut22_14), .ScanIn(nScanOut1487), .ScanOut(nScanOut1486), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1487 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_15), .NorthIn(nOut23_14), .SouthIn(nOut23_16), .EastIn(nOut24_15), .WestIn(nOut22_15), .ScanIn(nScanOut1488), .ScanOut(nScanOut1487), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1488 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_16), .NorthIn(nOut23_15), .SouthIn(nOut23_17), .EastIn(nOut24_16), .WestIn(nOut22_16), .ScanIn(nScanOut1489), .ScanOut(nScanOut1488), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1489 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_17), .NorthIn(nOut23_16), .SouthIn(nOut23_18), .EastIn(nOut24_17), .WestIn(nOut22_17), .ScanIn(nScanOut1490), .ScanOut(nScanOut1489), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1490 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_18), .NorthIn(nOut23_17), .SouthIn(nOut23_19), .EastIn(nOut24_18), .WestIn(nOut22_18), .ScanIn(nScanOut1491), .ScanOut(nScanOut1490), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1491 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_19), .NorthIn(nOut23_18), .SouthIn(nOut23_20), .EastIn(nOut24_19), .WestIn(nOut22_19), .ScanIn(nScanOut1492), .ScanOut(nScanOut1491), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1492 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_20), .NorthIn(nOut23_19), .SouthIn(nOut23_21), .EastIn(nOut24_20), .WestIn(nOut22_20), .ScanIn(nScanOut1493), .ScanOut(nScanOut1492), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1493 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_21), .NorthIn(nOut23_20), .SouthIn(nOut23_22), .EastIn(nOut24_21), .WestIn(nOut22_21), .ScanIn(nScanOut1494), .ScanOut(nScanOut1493), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1494 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_22), .NorthIn(nOut23_21), .SouthIn(nOut23_23), .EastIn(nOut24_22), .WestIn(nOut22_22), .ScanIn(nScanOut1495), .ScanOut(nScanOut1494), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1495 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_23), .NorthIn(nOut23_22), .SouthIn(nOut23_24), .EastIn(nOut24_23), .WestIn(nOut22_23), .ScanIn(nScanOut1496), .ScanOut(nScanOut1495), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1496 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_24), .NorthIn(nOut23_23), .SouthIn(nOut23_25), .EastIn(nOut24_24), .WestIn(nOut22_24), .ScanIn(nScanOut1497), .ScanOut(nScanOut1496), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1497 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_25), .NorthIn(nOut23_24), .SouthIn(nOut23_26), .EastIn(nOut24_25), .WestIn(nOut22_25), .ScanIn(nScanOut1498), .ScanOut(nScanOut1497), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1498 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_26), .NorthIn(nOut23_25), .SouthIn(nOut23_27), .EastIn(nOut24_26), .WestIn(nOut22_26), .ScanIn(nScanOut1499), .ScanOut(nScanOut1498), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1499 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_27), .NorthIn(nOut23_26), .SouthIn(nOut23_28), .EastIn(nOut24_27), .WestIn(nOut22_27), .ScanIn(nScanOut1500), .ScanOut(nScanOut1499), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1500 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_28), .NorthIn(nOut23_27), .SouthIn(nOut23_29), .EastIn(nOut24_28), .WestIn(nOut22_28), .ScanIn(nScanOut1501), .ScanOut(nScanOut1500), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1501 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_29), .NorthIn(nOut23_28), .SouthIn(nOut23_30), .EastIn(nOut24_29), .WestIn(nOut22_29), .ScanIn(nScanOut1502), .ScanOut(nScanOut1501), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1502 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_30), .NorthIn(nOut23_29), .SouthIn(nOut23_31), .EastIn(nOut24_30), .WestIn(nOut22_30), .ScanIn(nScanOut1503), .ScanOut(nScanOut1502), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1503 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_31), .NorthIn(nOut23_30), .SouthIn(nOut23_32), .EastIn(nOut24_31), .WestIn(nOut22_31), .ScanIn(nScanOut1504), .ScanOut(nScanOut1503), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1504 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_32), .NorthIn(nOut23_31), .SouthIn(nOut23_33), .EastIn(nOut24_32), .WestIn(nOut22_32), .ScanIn(nScanOut1505), .ScanOut(nScanOut1504), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1505 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_33), .NorthIn(nOut23_32), .SouthIn(nOut23_34), .EastIn(nOut24_33), .WestIn(nOut22_33), .ScanIn(nScanOut1506), .ScanOut(nScanOut1505), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1506 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_34), .NorthIn(nOut23_33), .SouthIn(nOut23_35), .EastIn(nOut24_34), .WestIn(nOut22_34), .ScanIn(nScanOut1507), .ScanOut(nScanOut1506), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1507 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_35), .NorthIn(nOut23_34), .SouthIn(nOut23_36), .EastIn(nOut24_35), .WestIn(nOut22_35), .ScanIn(nScanOut1508), .ScanOut(nScanOut1507), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1508 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_36), .NorthIn(nOut23_35), .SouthIn(nOut23_37), .EastIn(nOut24_36), .WestIn(nOut22_36), .ScanIn(nScanOut1509), .ScanOut(nScanOut1508), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1509 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_37), .NorthIn(nOut23_36), .SouthIn(nOut23_38), .EastIn(nOut24_37), .WestIn(nOut22_37), .ScanIn(nScanOut1510), .ScanOut(nScanOut1509), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1510 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_38), .NorthIn(nOut23_37), .SouthIn(nOut23_39), .EastIn(nOut24_38), .WestIn(nOut22_38), .ScanIn(nScanOut1511), .ScanOut(nScanOut1510), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1511 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_39), .NorthIn(nOut23_38), .SouthIn(nOut23_40), .EastIn(nOut24_39), .WestIn(nOut22_39), .ScanIn(nScanOut1512), .ScanOut(nScanOut1511), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1512 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_40), .NorthIn(nOut23_39), .SouthIn(nOut23_41), .EastIn(nOut24_40), .WestIn(nOut22_40), .ScanIn(nScanOut1513), .ScanOut(nScanOut1512), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1513 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_41), .NorthIn(nOut23_40), .SouthIn(nOut23_42), .EastIn(nOut24_41), .WestIn(nOut22_41), .ScanIn(nScanOut1514), .ScanOut(nScanOut1513), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1514 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_42), .NorthIn(nOut23_41), .SouthIn(nOut23_43), .EastIn(nOut24_42), .WestIn(nOut22_42), .ScanIn(nScanOut1515), .ScanOut(nScanOut1514), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1515 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_43), .NorthIn(nOut23_42), .SouthIn(nOut23_44), .EastIn(nOut24_43), .WestIn(nOut22_43), .ScanIn(nScanOut1516), .ScanOut(nScanOut1515), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1516 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_44), .NorthIn(nOut23_43), .SouthIn(nOut23_45), .EastIn(nOut24_44), .WestIn(nOut22_44), .ScanIn(nScanOut1517), .ScanOut(nScanOut1516), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1517 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_45), .NorthIn(nOut23_44), .SouthIn(nOut23_46), .EastIn(nOut24_45), .WestIn(nOut22_45), .ScanIn(nScanOut1518), .ScanOut(nScanOut1517), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1518 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_46), .NorthIn(nOut23_45), .SouthIn(nOut23_47), .EastIn(nOut24_46), .WestIn(nOut22_46), .ScanIn(nScanOut1519), .ScanOut(nScanOut1518), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1519 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_47), .NorthIn(nOut23_46), .SouthIn(nOut23_48), .EastIn(nOut24_47), .WestIn(nOut22_47), .ScanIn(nScanOut1520), .ScanOut(nScanOut1519), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1520 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_48), .NorthIn(nOut23_47), .SouthIn(nOut23_49), .EastIn(nOut24_48), .WestIn(nOut22_48), .ScanIn(nScanOut1521), .ScanOut(nScanOut1520), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1521 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_49), .NorthIn(nOut23_48), .SouthIn(nOut23_50), .EastIn(nOut24_49), .WestIn(nOut22_49), .ScanIn(nScanOut1522), .ScanOut(nScanOut1521), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1522 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_50), .NorthIn(nOut23_49), .SouthIn(nOut23_51), .EastIn(nOut24_50), .WestIn(nOut22_50), .ScanIn(nScanOut1523), .ScanOut(nScanOut1522), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1523 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_51), .NorthIn(nOut23_50), .SouthIn(nOut23_52), .EastIn(nOut24_51), .WestIn(nOut22_51), .ScanIn(nScanOut1524), .ScanOut(nScanOut1523), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1524 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_52), .NorthIn(nOut23_51), .SouthIn(nOut23_53), .EastIn(nOut24_52), .WestIn(nOut22_52), .ScanIn(nScanOut1525), .ScanOut(nScanOut1524), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1525 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_53), .NorthIn(nOut23_52), .SouthIn(nOut23_54), .EastIn(nOut24_53), .WestIn(nOut22_53), .ScanIn(nScanOut1526), .ScanOut(nScanOut1525), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1526 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_54), .NorthIn(nOut23_53), .SouthIn(nOut23_55), .EastIn(nOut24_54), .WestIn(nOut22_54), .ScanIn(nScanOut1527), .ScanOut(nScanOut1526), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1527 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_55), .NorthIn(nOut23_54), .SouthIn(nOut23_56), .EastIn(nOut24_55), .WestIn(nOut22_55), .ScanIn(nScanOut1528), .ScanOut(nScanOut1527), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1528 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_56), .NorthIn(nOut23_55), .SouthIn(nOut23_57), .EastIn(nOut24_56), .WestIn(nOut22_56), .ScanIn(nScanOut1529), .ScanOut(nScanOut1528), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1529 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_57), .NorthIn(nOut23_56), .SouthIn(nOut23_58), .EastIn(nOut24_57), .WestIn(nOut22_57), .ScanIn(nScanOut1530), .ScanOut(nScanOut1529), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1530 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_58), .NorthIn(nOut23_57), .SouthIn(nOut23_59), .EastIn(nOut24_58), .WestIn(nOut22_58), .ScanIn(nScanOut1531), .ScanOut(nScanOut1530), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1531 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_59), .NorthIn(nOut23_58), .SouthIn(nOut23_60), .EastIn(nOut24_59), .WestIn(nOut22_59), .ScanIn(nScanOut1532), .ScanOut(nScanOut1531), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1532 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_60), .NorthIn(nOut23_59), .SouthIn(nOut23_61), .EastIn(nOut24_60), .WestIn(nOut22_60), .ScanIn(nScanOut1533), .ScanOut(nScanOut1532), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1533 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_61), .NorthIn(nOut23_60), .SouthIn(nOut23_62), .EastIn(nOut24_61), .WestIn(nOut22_61), .ScanIn(nScanOut1534), .ScanOut(nScanOut1533), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1534 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut23_62), .NorthIn(nOut23_61), .SouthIn(nOut23_63), .EastIn(nOut24_62), .WestIn(nOut22_62), .ScanIn(nScanOut1535), .ScanOut(nScanOut1534), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1535 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut23_63), .ScanIn(nScanOut1536), .ScanOut(nScanOut1535), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1536 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut24_0), .ScanIn(nScanOut1537), .ScanOut(nScanOut1536), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1537 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_1), .NorthIn(nOut24_0), .SouthIn(nOut24_2), .EastIn(nOut25_1), .WestIn(nOut23_1), .ScanIn(nScanOut1538), .ScanOut(nScanOut1537), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1538 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_2), .NorthIn(nOut24_1), .SouthIn(nOut24_3), .EastIn(nOut25_2), .WestIn(nOut23_2), .ScanIn(nScanOut1539), .ScanOut(nScanOut1538), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1539 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_3), .NorthIn(nOut24_2), .SouthIn(nOut24_4), .EastIn(nOut25_3), .WestIn(nOut23_3), .ScanIn(nScanOut1540), .ScanOut(nScanOut1539), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1540 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_4), .NorthIn(nOut24_3), .SouthIn(nOut24_5), .EastIn(nOut25_4), .WestIn(nOut23_4), .ScanIn(nScanOut1541), .ScanOut(nScanOut1540), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1541 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_5), .NorthIn(nOut24_4), .SouthIn(nOut24_6), .EastIn(nOut25_5), .WestIn(nOut23_5), .ScanIn(nScanOut1542), .ScanOut(nScanOut1541), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1542 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_6), .NorthIn(nOut24_5), .SouthIn(nOut24_7), .EastIn(nOut25_6), .WestIn(nOut23_6), .ScanIn(nScanOut1543), .ScanOut(nScanOut1542), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1543 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_7), .NorthIn(nOut24_6), .SouthIn(nOut24_8), .EastIn(nOut25_7), .WestIn(nOut23_7), .ScanIn(nScanOut1544), .ScanOut(nScanOut1543), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1544 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_8), .NorthIn(nOut24_7), .SouthIn(nOut24_9), .EastIn(nOut25_8), .WestIn(nOut23_8), .ScanIn(nScanOut1545), .ScanOut(nScanOut1544), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1545 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_9), .NorthIn(nOut24_8), .SouthIn(nOut24_10), .EastIn(nOut25_9), .WestIn(nOut23_9), .ScanIn(nScanOut1546), .ScanOut(nScanOut1545), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1546 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_10), .NorthIn(nOut24_9), .SouthIn(nOut24_11), .EastIn(nOut25_10), .WestIn(nOut23_10), .ScanIn(nScanOut1547), .ScanOut(nScanOut1546), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1547 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_11), .NorthIn(nOut24_10), .SouthIn(nOut24_12), .EastIn(nOut25_11), .WestIn(nOut23_11), .ScanIn(nScanOut1548), .ScanOut(nScanOut1547), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1548 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_12), .NorthIn(nOut24_11), .SouthIn(nOut24_13), .EastIn(nOut25_12), .WestIn(nOut23_12), .ScanIn(nScanOut1549), .ScanOut(nScanOut1548), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1549 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_13), .NorthIn(nOut24_12), .SouthIn(nOut24_14), .EastIn(nOut25_13), .WestIn(nOut23_13), .ScanIn(nScanOut1550), .ScanOut(nScanOut1549), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1550 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_14), .NorthIn(nOut24_13), .SouthIn(nOut24_15), .EastIn(nOut25_14), .WestIn(nOut23_14), .ScanIn(nScanOut1551), .ScanOut(nScanOut1550), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1551 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_15), .NorthIn(nOut24_14), .SouthIn(nOut24_16), .EastIn(nOut25_15), .WestIn(nOut23_15), .ScanIn(nScanOut1552), .ScanOut(nScanOut1551), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1552 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_16), .NorthIn(nOut24_15), .SouthIn(nOut24_17), .EastIn(nOut25_16), .WestIn(nOut23_16), .ScanIn(nScanOut1553), .ScanOut(nScanOut1552), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1553 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_17), .NorthIn(nOut24_16), .SouthIn(nOut24_18), .EastIn(nOut25_17), .WestIn(nOut23_17), .ScanIn(nScanOut1554), .ScanOut(nScanOut1553), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1554 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_18), .NorthIn(nOut24_17), .SouthIn(nOut24_19), .EastIn(nOut25_18), .WestIn(nOut23_18), .ScanIn(nScanOut1555), .ScanOut(nScanOut1554), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1555 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_19), .NorthIn(nOut24_18), .SouthIn(nOut24_20), .EastIn(nOut25_19), .WestIn(nOut23_19), .ScanIn(nScanOut1556), .ScanOut(nScanOut1555), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1556 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_20), .NorthIn(nOut24_19), .SouthIn(nOut24_21), .EastIn(nOut25_20), .WestIn(nOut23_20), .ScanIn(nScanOut1557), .ScanOut(nScanOut1556), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1557 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_21), .NorthIn(nOut24_20), .SouthIn(nOut24_22), .EastIn(nOut25_21), .WestIn(nOut23_21), .ScanIn(nScanOut1558), .ScanOut(nScanOut1557), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1558 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_22), .NorthIn(nOut24_21), .SouthIn(nOut24_23), .EastIn(nOut25_22), .WestIn(nOut23_22), .ScanIn(nScanOut1559), .ScanOut(nScanOut1558), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1559 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_23), .NorthIn(nOut24_22), .SouthIn(nOut24_24), .EastIn(nOut25_23), .WestIn(nOut23_23), .ScanIn(nScanOut1560), .ScanOut(nScanOut1559), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1560 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_24), .NorthIn(nOut24_23), .SouthIn(nOut24_25), .EastIn(nOut25_24), .WestIn(nOut23_24), .ScanIn(nScanOut1561), .ScanOut(nScanOut1560), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1561 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_25), .NorthIn(nOut24_24), .SouthIn(nOut24_26), .EastIn(nOut25_25), .WestIn(nOut23_25), .ScanIn(nScanOut1562), .ScanOut(nScanOut1561), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1562 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_26), .NorthIn(nOut24_25), .SouthIn(nOut24_27), .EastIn(nOut25_26), .WestIn(nOut23_26), .ScanIn(nScanOut1563), .ScanOut(nScanOut1562), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1563 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_27), .NorthIn(nOut24_26), .SouthIn(nOut24_28), .EastIn(nOut25_27), .WestIn(nOut23_27), .ScanIn(nScanOut1564), .ScanOut(nScanOut1563), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1564 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_28), .NorthIn(nOut24_27), .SouthIn(nOut24_29), .EastIn(nOut25_28), .WestIn(nOut23_28), .ScanIn(nScanOut1565), .ScanOut(nScanOut1564), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1565 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_29), .NorthIn(nOut24_28), .SouthIn(nOut24_30), .EastIn(nOut25_29), .WestIn(nOut23_29), .ScanIn(nScanOut1566), .ScanOut(nScanOut1565), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1566 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_30), .NorthIn(nOut24_29), .SouthIn(nOut24_31), .EastIn(nOut25_30), .WestIn(nOut23_30), .ScanIn(nScanOut1567), .ScanOut(nScanOut1566), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1567 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_31), .NorthIn(nOut24_30), .SouthIn(nOut24_32), .EastIn(nOut25_31), .WestIn(nOut23_31), .ScanIn(nScanOut1568), .ScanOut(nScanOut1567), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1568 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_32), .NorthIn(nOut24_31), .SouthIn(nOut24_33), .EastIn(nOut25_32), .WestIn(nOut23_32), .ScanIn(nScanOut1569), .ScanOut(nScanOut1568), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1569 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_33), .NorthIn(nOut24_32), .SouthIn(nOut24_34), .EastIn(nOut25_33), .WestIn(nOut23_33), .ScanIn(nScanOut1570), .ScanOut(nScanOut1569), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1570 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_34), .NorthIn(nOut24_33), .SouthIn(nOut24_35), .EastIn(nOut25_34), .WestIn(nOut23_34), .ScanIn(nScanOut1571), .ScanOut(nScanOut1570), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1571 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_35), .NorthIn(nOut24_34), .SouthIn(nOut24_36), .EastIn(nOut25_35), .WestIn(nOut23_35), .ScanIn(nScanOut1572), .ScanOut(nScanOut1571), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1572 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_36), .NorthIn(nOut24_35), .SouthIn(nOut24_37), .EastIn(nOut25_36), .WestIn(nOut23_36), .ScanIn(nScanOut1573), .ScanOut(nScanOut1572), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1573 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_37), .NorthIn(nOut24_36), .SouthIn(nOut24_38), .EastIn(nOut25_37), .WestIn(nOut23_37), .ScanIn(nScanOut1574), .ScanOut(nScanOut1573), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1574 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_38), .NorthIn(nOut24_37), .SouthIn(nOut24_39), .EastIn(nOut25_38), .WestIn(nOut23_38), .ScanIn(nScanOut1575), .ScanOut(nScanOut1574), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1575 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_39), .NorthIn(nOut24_38), .SouthIn(nOut24_40), .EastIn(nOut25_39), .WestIn(nOut23_39), .ScanIn(nScanOut1576), .ScanOut(nScanOut1575), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1576 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_40), .NorthIn(nOut24_39), .SouthIn(nOut24_41), .EastIn(nOut25_40), .WestIn(nOut23_40), .ScanIn(nScanOut1577), .ScanOut(nScanOut1576), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1577 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_41), .NorthIn(nOut24_40), .SouthIn(nOut24_42), .EastIn(nOut25_41), .WestIn(nOut23_41), .ScanIn(nScanOut1578), .ScanOut(nScanOut1577), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1578 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_42), .NorthIn(nOut24_41), .SouthIn(nOut24_43), .EastIn(nOut25_42), .WestIn(nOut23_42), .ScanIn(nScanOut1579), .ScanOut(nScanOut1578), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1579 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_43), .NorthIn(nOut24_42), .SouthIn(nOut24_44), .EastIn(nOut25_43), .WestIn(nOut23_43), .ScanIn(nScanOut1580), .ScanOut(nScanOut1579), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1580 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_44), .NorthIn(nOut24_43), .SouthIn(nOut24_45), .EastIn(nOut25_44), .WestIn(nOut23_44), .ScanIn(nScanOut1581), .ScanOut(nScanOut1580), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1581 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_45), .NorthIn(nOut24_44), .SouthIn(nOut24_46), .EastIn(nOut25_45), .WestIn(nOut23_45), .ScanIn(nScanOut1582), .ScanOut(nScanOut1581), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1582 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_46), .NorthIn(nOut24_45), .SouthIn(nOut24_47), .EastIn(nOut25_46), .WestIn(nOut23_46), .ScanIn(nScanOut1583), .ScanOut(nScanOut1582), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1583 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_47), .NorthIn(nOut24_46), .SouthIn(nOut24_48), .EastIn(nOut25_47), .WestIn(nOut23_47), .ScanIn(nScanOut1584), .ScanOut(nScanOut1583), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1584 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_48), .NorthIn(nOut24_47), .SouthIn(nOut24_49), .EastIn(nOut25_48), .WestIn(nOut23_48), .ScanIn(nScanOut1585), .ScanOut(nScanOut1584), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1585 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_49), .NorthIn(nOut24_48), .SouthIn(nOut24_50), .EastIn(nOut25_49), .WestIn(nOut23_49), .ScanIn(nScanOut1586), .ScanOut(nScanOut1585), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1586 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_50), .NorthIn(nOut24_49), .SouthIn(nOut24_51), .EastIn(nOut25_50), .WestIn(nOut23_50), .ScanIn(nScanOut1587), .ScanOut(nScanOut1586), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1587 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_51), .NorthIn(nOut24_50), .SouthIn(nOut24_52), .EastIn(nOut25_51), .WestIn(nOut23_51), .ScanIn(nScanOut1588), .ScanOut(nScanOut1587), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1588 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_52), .NorthIn(nOut24_51), .SouthIn(nOut24_53), .EastIn(nOut25_52), .WestIn(nOut23_52), .ScanIn(nScanOut1589), .ScanOut(nScanOut1588), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1589 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_53), .NorthIn(nOut24_52), .SouthIn(nOut24_54), .EastIn(nOut25_53), .WestIn(nOut23_53), .ScanIn(nScanOut1590), .ScanOut(nScanOut1589), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1590 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_54), .NorthIn(nOut24_53), .SouthIn(nOut24_55), .EastIn(nOut25_54), .WestIn(nOut23_54), .ScanIn(nScanOut1591), .ScanOut(nScanOut1590), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1591 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_55), .NorthIn(nOut24_54), .SouthIn(nOut24_56), .EastIn(nOut25_55), .WestIn(nOut23_55), .ScanIn(nScanOut1592), .ScanOut(nScanOut1591), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1592 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_56), .NorthIn(nOut24_55), .SouthIn(nOut24_57), .EastIn(nOut25_56), .WestIn(nOut23_56), .ScanIn(nScanOut1593), .ScanOut(nScanOut1592), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1593 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_57), .NorthIn(nOut24_56), .SouthIn(nOut24_58), .EastIn(nOut25_57), .WestIn(nOut23_57), .ScanIn(nScanOut1594), .ScanOut(nScanOut1593), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1594 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_58), .NorthIn(nOut24_57), .SouthIn(nOut24_59), .EastIn(nOut25_58), .WestIn(nOut23_58), .ScanIn(nScanOut1595), .ScanOut(nScanOut1594), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1595 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_59), .NorthIn(nOut24_58), .SouthIn(nOut24_60), .EastIn(nOut25_59), .WestIn(nOut23_59), .ScanIn(nScanOut1596), .ScanOut(nScanOut1595), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1596 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_60), .NorthIn(nOut24_59), .SouthIn(nOut24_61), .EastIn(nOut25_60), .WestIn(nOut23_60), .ScanIn(nScanOut1597), .ScanOut(nScanOut1596), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1597 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_61), .NorthIn(nOut24_60), .SouthIn(nOut24_62), .EastIn(nOut25_61), .WestIn(nOut23_61), .ScanIn(nScanOut1598), .ScanOut(nScanOut1597), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1598 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut24_62), .NorthIn(nOut24_61), .SouthIn(nOut24_63), .EastIn(nOut25_62), .WestIn(nOut23_62), .ScanIn(nScanOut1599), .ScanOut(nScanOut1598), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1599 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut24_63), .ScanIn(nScanOut1600), .ScanOut(nScanOut1599), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1600 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut25_0), .ScanIn(nScanOut1601), .ScanOut(nScanOut1600), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1601 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_1), .NorthIn(nOut25_0), .SouthIn(nOut25_2), .EastIn(nOut26_1), .WestIn(nOut24_1), .ScanIn(nScanOut1602), .ScanOut(nScanOut1601), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1602 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_2), .NorthIn(nOut25_1), .SouthIn(nOut25_3), .EastIn(nOut26_2), .WestIn(nOut24_2), .ScanIn(nScanOut1603), .ScanOut(nScanOut1602), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1603 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_3), .NorthIn(nOut25_2), .SouthIn(nOut25_4), .EastIn(nOut26_3), .WestIn(nOut24_3), .ScanIn(nScanOut1604), .ScanOut(nScanOut1603), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1604 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_4), .NorthIn(nOut25_3), .SouthIn(nOut25_5), .EastIn(nOut26_4), .WestIn(nOut24_4), .ScanIn(nScanOut1605), .ScanOut(nScanOut1604), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1605 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_5), .NorthIn(nOut25_4), .SouthIn(nOut25_6), .EastIn(nOut26_5), .WestIn(nOut24_5), .ScanIn(nScanOut1606), .ScanOut(nScanOut1605), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1606 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_6), .NorthIn(nOut25_5), .SouthIn(nOut25_7), .EastIn(nOut26_6), .WestIn(nOut24_6), .ScanIn(nScanOut1607), .ScanOut(nScanOut1606), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1607 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_7), .NorthIn(nOut25_6), .SouthIn(nOut25_8), .EastIn(nOut26_7), .WestIn(nOut24_7), .ScanIn(nScanOut1608), .ScanOut(nScanOut1607), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1608 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_8), .NorthIn(nOut25_7), .SouthIn(nOut25_9), .EastIn(nOut26_8), .WestIn(nOut24_8), .ScanIn(nScanOut1609), .ScanOut(nScanOut1608), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1609 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_9), .NorthIn(nOut25_8), .SouthIn(nOut25_10), .EastIn(nOut26_9), .WestIn(nOut24_9), .ScanIn(nScanOut1610), .ScanOut(nScanOut1609), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1610 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_10), .NorthIn(nOut25_9), .SouthIn(nOut25_11), .EastIn(nOut26_10), .WestIn(nOut24_10), .ScanIn(nScanOut1611), .ScanOut(nScanOut1610), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1611 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_11), .NorthIn(nOut25_10), .SouthIn(nOut25_12), .EastIn(nOut26_11), .WestIn(nOut24_11), .ScanIn(nScanOut1612), .ScanOut(nScanOut1611), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1612 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_12), .NorthIn(nOut25_11), .SouthIn(nOut25_13), .EastIn(nOut26_12), .WestIn(nOut24_12), .ScanIn(nScanOut1613), .ScanOut(nScanOut1612), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1613 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_13), .NorthIn(nOut25_12), .SouthIn(nOut25_14), .EastIn(nOut26_13), .WestIn(nOut24_13), .ScanIn(nScanOut1614), .ScanOut(nScanOut1613), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1614 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_14), .NorthIn(nOut25_13), .SouthIn(nOut25_15), .EastIn(nOut26_14), .WestIn(nOut24_14), .ScanIn(nScanOut1615), .ScanOut(nScanOut1614), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1615 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_15), .NorthIn(nOut25_14), .SouthIn(nOut25_16), .EastIn(nOut26_15), .WestIn(nOut24_15), .ScanIn(nScanOut1616), .ScanOut(nScanOut1615), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1616 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_16), .NorthIn(nOut25_15), .SouthIn(nOut25_17), .EastIn(nOut26_16), .WestIn(nOut24_16), .ScanIn(nScanOut1617), .ScanOut(nScanOut1616), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1617 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_17), .NorthIn(nOut25_16), .SouthIn(nOut25_18), .EastIn(nOut26_17), .WestIn(nOut24_17), .ScanIn(nScanOut1618), .ScanOut(nScanOut1617), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1618 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_18), .NorthIn(nOut25_17), .SouthIn(nOut25_19), .EastIn(nOut26_18), .WestIn(nOut24_18), .ScanIn(nScanOut1619), .ScanOut(nScanOut1618), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1619 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_19), .NorthIn(nOut25_18), .SouthIn(nOut25_20), .EastIn(nOut26_19), .WestIn(nOut24_19), .ScanIn(nScanOut1620), .ScanOut(nScanOut1619), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1620 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_20), .NorthIn(nOut25_19), .SouthIn(nOut25_21), .EastIn(nOut26_20), .WestIn(nOut24_20), .ScanIn(nScanOut1621), .ScanOut(nScanOut1620), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1621 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_21), .NorthIn(nOut25_20), .SouthIn(nOut25_22), .EastIn(nOut26_21), .WestIn(nOut24_21), .ScanIn(nScanOut1622), .ScanOut(nScanOut1621), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1622 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_22), .NorthIn(nOut25_21), .SouthIn(nOut25_23), .EastIn(nOut26_22), .WestIn(nOut24_22), .ScanIn(nScanOut1623), .ScanOut(nScanOut1622), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1623 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_23), .NorthIn(nOut25_22), .SouthIn(nOut25_24), .EastIn(nOut26_23), .WestIn(nOut24_23), .ScanIn(nScanOut1624), .ScanOut(nScanOut1623), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1624 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_24), .NorthIn(nOut25_23), .SouthIn(nOut25_25), .EastIn(nOut26_24), .WestIn(nOut24_24), .ScanIn(nScanOut1625), .ScanOut(nScanOut1624), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1625 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_25), .NorthIn(nOut25_24), .SouthIn(nOut25_26), .EastIn(nOut26_25), .WestIn(nOut24_25), .ScanIn(nScanOut1626), .ScanOut(nScanOut1625), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1626 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_26), .NorthIn(nOut25_25), .SouthIn(nOut25_27), .EastIn(nOut26_26), .WestIn(nOut24_26), .ScanIn(nScanOut1627), .ScanOut(nScanOut1626), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1627 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_27), .NorthIn(nOut25_26), .SouthIn(nOut25_28), .EastIn(nOut26_27), .WestIn(nOut24_27), .ScanIn(nScanOut1628), .ScanOut(nScanOut1627), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1628 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_28), .NorthIn(nOut25_27), .SouthIn(nOut25_29), .EastIn(nOut26_28), .WestIn(nOut24_28), .ScanIn(nScanOut1629), .ScanOut(nScanOut1628), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1629 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_29), .NorthIn(nOut25_28), .SouthIn(nOut25_30), .EastIn(nOut26_29), .WestIn(nOut24_29), .ScanIn(nScanOut1630), .ScanOut(nScanOut1629), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1630 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_30), .NorthIn(nOut25_29), .SouthIn(nOut25_31), .EastIn(nOut26_30), .WestIn(nOut24_30), .ScanIn(nScanOut1631), .ScanOut(nScanOut1630), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1631 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_31), .NorthIn(nOut25_30), .SouthIn(nOut25_32), .EastIn(nOut26_31), .WestIn(nOut24_31), .ScanIn(nScanOut1632), .ScanOut(nScanOut1631), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1632 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_32), .NorthIn(nOut25_31), .SouthIn(nOut25_33), .EastIn(nOut26_32), .WestIn(nOut24_32), .ScanIn(nScanOut1633), .ScanOut(nScanOut1632), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1633 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_33), .NorthIn(nOut25_32), .SouthIn(nOut25_34), .EastIn(nOut26_33), .WestIn(nOut24_33), .ScanIn(nScanOut1634), .ScanOut(nScanOut1633), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1634 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_34), .NorthIn(nOut25_33), .SouthIn(nOut25_35), .EastIn(nOut26_34), .WestIn(nOut24_34), .ScanIn(nScanOut1635), .ScanOut(nScanOut1634), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1635 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_35), .NorthIn(nOut25_34), .SouthIn(nOut25_36), .EastIn(nOut26_35), .WestIn(nOut24_35), .ScanIn(nScanOut1636), .ScanOut(nScanOut1635), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1636 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_36), .NorthIn(nOut25_35), .SouthIn(nOut25_37), .EastIn(nOut26_36), .WestIn(nOut24_36), .ScanIn(nScanOut1637), .ScanOut(nScanOut1636), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1637 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_37), .NorthIn(nOut25_36), .SouthIn(nOut25_38), .EastIn(nOut26_37), .WestIn(nOut24_37), .ScanIn(nScanOut1638), .ScanOut(nScanOut1637), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1638 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_38), .NorthIn(nOut25_37), .SouthIn(nOut25_39), .EastIn(nOut26_38), .WestIn(nOut24_38), .ScanIn(nScanOut1639), .ScanOut(nScanOut1638), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1639 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_39), .NorthIn(nOut25_38), .SouthIn(nOut25_40), .EastIn(nOut26_39), .WestIn(nOut24_39), .ScanIn(nScanOut1640), .ScanOut(nScanOut1639), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1640 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_40), .NorthIn(nOut25_39), .SouthIn(nOut25_41), .EastIn(nOut26_40), .WestIn(nOut24_40), .ScanIn(nScanOut1641), .ScanOut(nScanOut1640), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1641 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_41), .NorthIn(nOut25_40), .SouthIn(nOut25_42), .EastIn(nOut26_41), .WestIn(nOut24_41), .ScanIn(nScanOut1642), .ScanOut(nScanOut1641), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1642 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_42), .NorthIn(nOut25_41), .SouthIn(nOut25_43), .EastIn(nOut26_42), .WestIn(nOut24_42), .ScanIn(nScanOut1643), .ScanOut(nScanOut1642), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1643 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_43), .NorthIn(nOut25_42), .SouthIn(nOut25_44), .EastIn(nOut26_43), .WestIn(nOut24_43), .ScanIn(nScanOut1644), .ScanOut(nScanOut1643), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1644 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_44), .NorthIn(nOut25_43), .SouthIn(nOut25_45), .EastIn(nOut26_44), .WestIn(nOut24_44), .ScanIn(nScanOut1645), .ScanOut(nScanOut1644), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1645 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_45), .NorthIn(nOut25_44), .SouthIn(nOut25_46), .EastIn(nOut26_45), .WestIn(nOut24_45), .ScanIn(nScanOut1646), .ScanOut(nScanOut1645), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1646 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_46), .NorthIn(nOut25_45), .SouthIn(nOut25_47), .EastIn(nOut26_46), .WestIn(nOut24_46), .ScanIn(nScanOut1647), .ScanOut(nScanOut1646), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1647 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_47), .NorthIn(nOut25_46), .SouthIn(nOut25_48), .EastIn(nOut26_47), .WestIn(nOut24_47), .ScanIn(nScanOut1648), .ScanOut(nScanOut1647), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1648 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_48), .NorthIn(nOut25_47), .SouthIn(nOut25_49), .EastIn(nOut26_48), .WestIn(nOut24_48), .ScanIn(nScanOut1649), .ScanOut(nScanOut1648), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1649 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_49), .NorthIn(nOut25_48), .SouthIn(nOut25_50), .EastIn(nOut26_49), .WestIn(nOut24_49), .ScanIn(nScanOut1650), .ScanOut(nScanOut1649), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1650 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_50), .NorthIn(nOut25_49), .SouthIn(nOut25_51), .EastIn(nOut26_50), .WestIn(nOut24_50), .ScanIn(nScanOut1651), .ScanOut(nScanOut1650), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1651 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_51), .NorthIn(nOut25_50), .SouthIn(nOut25_52), .EastIn(nOut26_51), .WestIn(nOut24_51), .ScanIn(nScanOut1652), .ScanOut(nScanOut1651), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1652 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_52), .NorthIn(nOut25_51), .SouthIn(nOut25_53), .EastIn(nOut26_52), .WestIn(nOut24_52), .ScanIn(nScanOut1653), .ScanOut(nScanOut1652), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1653 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_53), .NorthIn(nOut25_52), .SouthIn(nOut25_54), .EastIn(nOut26_53), .WestIn(nOut24_53), .ScanIn(nScanOut1654), .ScanOut(nScanOut1653), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1654 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_54), .NorthIn(nOut25_53), .SouthIn(nOut25_55), .EastIn(nOut26_54), .WestIn(nOut24_54), .ScanIn(nScanOut1655), .ScanOut(nScanOut1654), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1655 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_55), .NorthIn(nOut25_54), .SouthIn(nOut25_56), .EastIn(nOut26_55), .WestIn(nOut24_55), .ScanIn(nScanOut1656), .ScanOut(nScanOut1655), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1656 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_56), .NorthIn(nOut25_55), .SouthIn(nOut25_57), .EastIn(nOut26_56), .WestIn(nOut24_56), .ScanIn(nScanOut1657), .ScanOut(nScanOut1656), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1657 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_57), .NorthIn(nOut25_56), .SouthIn(nOut25_58), .EastIn(nOut26_57), .WestIn(nOut24_57), .ScanIn(nScanOut1658), .ScanOut(nScanOut1657), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1658 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_58), .NorthIn(nOut25_57), .SouthIn(nOut25_59), .EastIn(nOut26_58), .WestIn(nOut24_58), .ScanIn(nScanOut1659), .ScanOut(nScanOut1658), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1659 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_59), .NorthIn(nOut25_58), .SouthIn(nOut25_60), .EastIn(nOut26_59), .WestIn(nOut24_59), .ScanIn(nScanOut1660), .ScanOut(nScanOut1659), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1660 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_60), .NorthIn(nOut25_59), .SouthIn(nOut25_61), .EastIn(nOut26_60), .WestIn(nOut24_60), .ScanIn(nScanOut1661), .ScanOut(nScanOut1660), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1661 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_61), .NorthIn(nOut25_60), .SouthIn(nOut25_62), .EastIn(nOut26_61), .WestIn(nOut24_61), .ScanIn(nScanOut1662), .ScanOut(nScanOut1661), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1662 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut25_62), .NorthIn(nOut25_61), .SouthIn(nOut25_63), .EastIn(nOut26_62), .WestIn(nOut24_62), .ScanIn(nScanOut1663), .ScanOut(nScanOut1662), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1663 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut25_63), .ScanIn(nScanOut1664), .ScanOut(nScanOut1663), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1664 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut26_0), .ScanIn(nScanOut1665), .ScanOut(nScanOut1664), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1665 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_1), .NorthIn(nOut26_0), .SouthIn(nOut26_2), .EastIn(nOut27_1), .WestIn(nOut25_1), .ScanIn(nScanOut1666), .ScanOut(nScanOut1665), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1666 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_2), .NorthIn(nOut26_1), .SouthIn(nOut26_3), .EastIn(nOut27_2), .WestIn(nOut25_2), .ScanIn(nScanOut1667), .ScanOut(nScanOut1666), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1667 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_3), .NorthIn(nOut26_2), .SouthIn(nOut26_4), .EastIn(nOut27_3), .WestIn(nOut25_3), .ScanIn(nScanOut1668), .ScanOut(nScanOut1667), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1668 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_4), .NorthIn(nOut26_3), .SouthIn(nOut26_5), .EastIn(nOut27_4), .WestIn(nOut25_4), .ScanIn(nScanOut1669), .ScanOut(nScanOut1668), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1669 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_5), .NorthIn(nOut26_4), .SouthIn(nOut26_6), .EastIn(nOut27_5), .WestIn(nOut25_5), .ScanIn(nScanOut1670), .ScanOut(nScanOut1669), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1670 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_6), .NorthIn(nOut26_5), .SouthIn(nOut26_7), .EastIn(nOut27_6), .WestIn(nOut25_6), .ScanIn(nScanOut1671), .ScanOut(nScanOut1670), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1671 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_7), .NorthIn(nOut26_6), .SouthIn(nOut26_8), .EastIn(nOut27_7), .WestIn(nOut25_7), .ScanIn(nScanOut1672), .ScanOut(nScanOut1671), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1672 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_8), .NorthIn(nOut26_7), .SouthIn(nOut26_9), .EastIn(nOut27_8), .WestIn(nOut25_8), .ScanIn(nScanOut1673), .ScanOut(nScanOut1672), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1673 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_9), .NorthIn(nOut26_8), .SouthIn(nOut26_10), .EastIn(nOut27_9), .WestIn(nOut25_9), .ScanIn(nScanOut1674), .ScanOut(nScanOut1673), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1674 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_10), .NorthIn(nOut26_9), .SouthIn(nOut26_11), .EastIn(nOut27_10), .WestIn(nOut25_10), .ScanIn(nScanOut1675), .ScanOut(nScanOut1674), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1675 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_11), .NorthIn(nOut26_10), .SouthIn(nOut26_12), .EastIn(nOut27_11), .WestIn(nOut25_11), .ScanIn(nScanOut1676), .ScanOut(nScanOut1675), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1676 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_12), .NorthIn(nOut26_11), .SouthIn(nOut26_13), .EastIn(nOut27_12), .WestIn(nOut25_12), .ScanIn(nScanOut1677), .ScanOut(nScanOut1676), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1677 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_13), .NorthIn(nOut26_12), .SouthIn(nOut26_14), .EastIn(nOut27_13), .WestIn(nOut25_13), .ScanIn(nScanOut1678), .ScanOut(nScanOut1677), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1678 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_14), .NorthIn(nOut26_13), .SouthIn(nOut26_15), .EastIn(nOut27_14), .WestIn(nOut25_14), .ScanIn(nScanOut1679), .ScanOut(nScanOut1678), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1679 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_15), .NorthIn(nOut26_14), .SouthIn(nOut26_16), .EastIn(nOut27_15), .WestIn(nOut25_15), .ScanIn(nScanOut1680), .ScanOut(nScanOut1679), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1680 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_16), .NorthIn(nOut26_15), .SouthIn(nOut26_17), .EastIn(nOut27_16), .WestIn(nOut25_16), .ScanIn(nScanOut1681), .ScanOut(nScanOut1680), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1681 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_17), .NorthIn(nOut26_16), .SouthIn(nOut26_18), .EastIn(nOut27_17), .WestIn(nOut25_17), .ScanIn(nScanOut1682), .ScanOut(nScanOut1681), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1682 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_18), .NorthIn(nOut26_17), .SouthIn(nOut26_19), .EastIn(nOut27_18), .WestIn(nOut25_18), .ScanIn(nScanOut1683), .ScanOut(nScanOut1682), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1683 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_19), .NorthIn(nOut26_18), .SouthIn(nOut26_20), .EastIn(nOut27_19), .WestIn(nOut25_19), .ScanIn(nScanOut1684), .ScanOut(nScanOut1683), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1684 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_20), .NorthIn(nOut26_19), .SouthIn(nOut26_21), .EastIn(nOut27_20), .WestIn(nOut25_20), .ScanIn(nScanOut1685), .ScanOut(nScanOut1684), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1685 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_21), .NorthIn(nOut26_20), .SouthIn(nOut26_22), .EastIn(nOut27_21), .WestIn(nOut25_21), .ScanIn(nScanOut1686), .ScanOut(nScanOut1685), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1686 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_22), .NorthIn(nOut26_21), .SouthIn(nOut26_23), .EastIn(nOut27_22), .WestIn(nOut25_22), .ScanIn(nScanOut1687), .ScanOut(nScanOut1686), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1687 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_23), .NorthIn(nOut26_22), .SouthIn(nOut26_24), .EastIn(nOut27_23), .WestIn(nOut25_23), .ScanIn(nScanOut1688), .ScanOut(nScanOut1687), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1688 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_24), .NorthIn(nOut26_23), .SouthIn(nOut26_25), .EastIn(nOut27_24), .WestIn(nOut25_24), .ScanIn(nScanOut1689), .ScanOut(nScanOut1688), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1689 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_25), .NorthIn(nOut26_24), .SouthIn(nOut26_26), .EastIn(nOut27_25), .WestIn(nOut25_25), .ScanIn(nScanOut1690), .ScanOut(nScanOut1689), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1690 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_26), .NorthIn(nOut26_25), .SouthIn(nOut26_27), .EastIn(nOut27_26), .WestIn(nOut25_26), .ScanIn(nScanOut1691), .ScanOut(nScanOut1690), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1691 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_27), .NorthIn(nOut26_26), .SouthIn(nOut26_28), .EastIn(nOut27_27), .WestIn(nOut25_27), .ScanIn(nScanOut1692), .ScanOut(nScanOut1691), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1692 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_28), .NorthIn(nOut26_27), .SouthIn(nOut26_29), .EastIn(nOut27_28), .WestIn(nOut25_28), .ScanIn(nScanOut1693), .ScanOut(nScanOut1692), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1693 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_29), .NorthIn(nOut26_28), .SouthIn(nOut26_30), .EastIn(nOut27_29), .WestIn(nOut25_29), .ScanIn(nScanOut1694), .ScanOut(nScanOut1693), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1694 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_30), .NorthIn(nOut26_29), .SouthIn(nOut26_31), .EastIn(nOut27_30), .WestIn(nOut25_30), .ScanIn(nScanOut1695), .ScanOut(nScanOut1694), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1695 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_31), .NorthIn(nOut26_30), .SouthIn(nOut26_32), .EastIn(nOut27_31), .WestIn(nOut25_31), .ScanIn(nScanOut1696), .ScanOut(nScanOut1695), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1696 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_32), .NorthIn(nOut26_31), .SouthIn(nOut26_33), .EastIn(nOut27_32), .WestIn(nOut25_32), .ScanIn(nScanOut1697), .ScanOut(nScanOut1696), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1697 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_33), .NorthIn(nOut26_32), .SouthIn(nOut26_34), .EastIn(nOut27_33), .WestIn(nOut25_33), .ScanIn(nScanOut1698), .ScanOut(nScanOut1697), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1698 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_34), .NorthIn(nOut26_33), .SouthIn(nOut26_35), .EastIn(nOut27_34), .WestIn(nOut25_34), .ScanIn(nScanOut1699), .ScanOut(nScanOut1698), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1699 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_35), .NorthIn(nOut26_34), .SouthIn(nOut26_36), .EastIn(nOut27_35), .WestIn(nOut25_35), .ScanIn(nScanOut1700), .ScanOut(nScanOut1699), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1700 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_36), .NorthIn(nOut26_35), .SouthIn(nOut26_37), .EastIn(nOut27_36), .WestIn(nOut25_36), .ScanIn(nScanOut1701), .ScanOut(nScanOut1700), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1701 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_37), .NorthIn(nOut26_36), .SouthIn(nOut26_38), .EastIn(nOut27_37), .WestIn(nOut25_37), .ScanIn(nScanOut1702), .ScanOut(nScanOut1701), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1702 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_38), .NorthIn(nOut26_37), .SouthIn(nOut26_39), .EastIn(nOut27_38), .WestIn(nOut25_38), .ScanIn(nScanOut1703), .ScanOut(nScanOut1702), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1703 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_39), .NorthIn(nOut26_38), .SouthIn(nOut26_40), .EastIn(nOut27_39), .WestIn(nOut25_39), .ScanIn(nScanOut1704), .ScanOut(nScanOut1703), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1704 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_40), .NorthIn(nOut26_39), .SouthIn(nOut26_41), .EastIn(nOut27_40), .WestIn(nOut25_40), .ScanIn(nScanOut1705), .ScanOut(nScanOut1704), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1705 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_41), .NorthIn(nOut26_40), .SouthIn(nOut26_42), .EastIn(nOut27_41), .WestIn(nOut25_41), .ScanIn(nScanOut1706), .ScanOut(nScanOut1705), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1706 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_42), .NorthIn(nOut26_41), .SouthIn(nOut26_43), .EastIn(nOut27_42), .WestIn(nOut25_42), .ScanIn(nScanOut1707), .ScanOut(nScanOut1706), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1707 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_43), .NorthIn(nOut26_42), .SouthIn(nOut26_44), .EastIn(nOut27_43), .WestIn(nOut25_43), .ScanIn(nScanOut1708), .ScanOut(nScanOut1707), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1708 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_44), .NorthIn(nOut26_43), .SouthIn(nOut26_45), .EastIn(nOut27_44), .WestIn(nOut25_44), .ScanIn(nScanOut1709), .ScanOut(nScanOut1708), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1709 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_45), .NorthIn(nOut26_44), .SouthIn(nOut26_46), .EastIn(nOut27_45), .WestIn(nOut25_45), .ScanIn(nScanOut1710), .ScanOut(nScanOut1709), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1710 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_46), .NorthIn(nOut26_45), .SouthIn(nOut26_47), .EastIn(nOut27_46), .WestIn(nOut25_46), .ScanIn(nScanOut1711), .ScanOut(nScanOut1710), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1711 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_47), .NorthIn(nOut26_46), .SouthIn(nOut26_48), .EastIn(nOut27_47), .WestIn(nOut25_47), .ScanIn(nScanOut1712), .ScanOut(nScanOut1711), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1712 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_48), .NorthIn(nOut26_47), .SouthIn(nOut26_49), .EastIn(nOut27_48), .WestIn(nOut25_48), .ScanIn(nScanOut1713), .ScanOut(nScanOut1712), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1713 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_49), .NorthIn(nOut26_48), .SouthIn(nOut26_50), .EastIn(nOut27_49), .WestIn(nOut25_49), .ScanIn(nScanOut1714), .ScanOut(nScanOut1713), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1714 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_50), .NorthIn(nOut26_49), .SouthIn(nOut26_51), .EastIn(nOut27_50), .WestIn(nOut25_50), .ScanIn(nScanOut1715), .ScanOut(nScanOut1714), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1715 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_51), .NorthIn(nOut26_50), .SouthIn(nOut26_52), .EastIn(nOut27_51), .WestIn(nOut25_51), .ScanIn(nScanOut1716), .ScanOut(nScanOut1715), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1716 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_52), .NorthIn(nOut26_51), .SouthIn(nOut26_53), .EastIn(nOut27_52), .WestIn(nOut25_52), .ScanIn(nScanOut1717), .ScanOut(nScanOut1716), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1717 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_53), .NorthIn(nOut26_52), .SouthIn(nOut26_54), .EastIn(nOut27_53), .WestIn(nOut25_53), .ScanIn(nScanOut1718), .ScanOut(nScanOut1717), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1718 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_54), .NorthIn(nOut26_53), .SouthIn(nOut26_55), .EastIn(nOut27_54), .WestIn(nOut25_54), .ScanIn(nScanOut1719), .ScanOut(nScanOut1718), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1719 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_55), .NorthIn(nOut26_54), .SouthIn(nOut26_56), .EastIn(nOut27_55), .WestIn(nOut25_55), .ScanIn(nScanOut1720), .ScanOut(nScanOut1719), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1720 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_56), .NorthIn(nOut26_55), .SouthIn(nOut26_57), .EastIn(nOut27_56), .WestIn(nOut25_56), .ScanIn(nScanOut1721), .ScanOut(nScanOut1720), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1721 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_57), .NorthIn(nOut26_56), .SouthIn(nOut26_58), .EastIn(nOut27_57), .WestIn(nOut25_57), .ScanIn(nScanOut1722), .ScanOut(nScanOut1721), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1722 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_58), .NorthIn(nOut26_57), .SouthIn(nOut26_59), .EastIn(nOut27_58), .WestIn(nOut25_58), .ScanIn(nScanOut1723), .ScanOut(nScanOut1722), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1723 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_59), .NorthIn(nOut26_58), .SouthIn(nOut26_60), .EastIn(nOut27_59), .WestIn(nOut25_59), .ScanIn(nScanOut1724), .ScanOut(nScanOut1723), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1724 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_60), .NorthIn(nOut26_59), .SouthIn(nOut26_61), .EastIn(nOut27_60), .WestIn(nOut25_60), .ScanIn(nScanOut1725), .ScanOut(nScanOut1724), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1725 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_61), .NorthIn(nOut26_60), .SouthIn(nOut26_62), .EastIn(nOut27_61), .WestIn(nOut25_61), .ScanIn(nScanOut1726), .ScanOut(nScanOut1725), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1726 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut26_62), .NorthIn(nOut26_61), .SouthIn(nOut26_63), .EastIn(nOut27_62), .WestIn(nOut25_62), .ScanIn(nScanOut1727), .ScanOut(nScanOut1726), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1727 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut26_63), .ScanIn(nScanOut1728), .ScanOut(nScanOut1727), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1728 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut27_0), .ScanIn(nScanOut1729), .ScanOut(nScanOut1728), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1729 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_1), .NorthIn(nOut27_0), .SouthIn(nOut27_2), .EastIn(nOut28_1), .WestIn(nOut26_1), .ScanIn(nScanOut1730), .ScanOut(nScanOut1729), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1730 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_2), .NorthIn(nOut27_1), .SouthIn(nOut27_3), .EastIn(nOut28_2), .WestIn(nOut26_2), .ScanIn(nScanOut1731), .ScanOut(nScanOut1730), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1731 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_3), .NorthIn(nOut27_2), .SouthIn(nOut27_4), .EastIn(nOut28_3), .WestIn(nOut26_3), .ScanIn(nScanOut1732), .ScanOut(nScanOut1731), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1732 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_4), .NorthIn(nOut27_3), .SouthIn(nOut27_5), .EastIn(nOut28_4), .WestIn(nOut26_4), .ScanIn(nScanOut1733), .ScanOut(nScanOut1732), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1733 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_5), .NorthIn(nOut27_4), .SouthIn(nOut27_6), .EastIn(nOut28_5), .WestIn(nOut26_5), .ScanIn(nScanOut1734), .ScanOut(nScanOut1733), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1734 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_6), .NorthIn(nOut27_5), .SouthIn(nOut27_7), .EastIn(nOut28_6), .WestIn(nOut26_6), .ScanIn(nScanOut1735), .ScanOut(nScanOut1734), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1735 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_7), .NorthIn(nOut27_6), .SouthIn(nOut27_8), .EastIn(nOut28_7), .WestIn(nOut26_7), .ScanIn(nScanOut1736), .ScanOut(nScanOut1735), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1736 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_8), .NorthIn(nOut27_7), .SouthIn(nOut27_9), .EastIn(nOut28_8), .WestIn(nOut26_8), .ScanIn(nScanOut1737), .ScanOut(nScanOut1736), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1737 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_9), .NorthIn(nOut27_8), .SouthIn(nOut27_10), .EastIn(nOut28_9), .WestIn(nOut26_9), .ScanIn(nScanOut1738), .ScanOut(nScanOut1737), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1738 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_10), .NorthIn(nOut27_9), .SouthIn(nOut27_11), .EastIn(nOut28_10), .WestIn(nOut26_10), .ScanIn(nScanOut1739), .ScanOut(nScanOut1738), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1739 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_11), .NorthIn(nOut27_10), .SouthIn(nOut27_12), .EastIn(nOut28_11), .WestIn(nOut26_11), .ScanIn(nScanOut1740), .ScanOut(nScanOut1739), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1740 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_12), .NorthIn(nOut27_11), .SouthIn(nOut27_13), .EastIn(nOut28_12), .WestIn(nOut26_12), .ScanIn(nScanOut1741), .ScanOut(nScanOut1740), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1741 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_13), .NorthIn(nOut27_12), .SouthIn(nOut27_14), .EastIn(nOut28_13), .WestIn(nOut26_13), .ScanIn(nScanOut1742), .ScanOut(nScanOut1741), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1742 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_14), .NorthIn(nOut27_13), .SouthIn(nOut27_15), .EastIn(nOut28_14), .WestIn(nOut26_14), .ScanIn(nScanOut1743), .ScanOut(nScanOut1742), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1743 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_15), .NorthIn(nOut27_14), .SouthIn(nOut27_16), .EastIn(nOut28_15), .WestIn(nOut26_15), .ScanIn(nScanOut1744), .ScanOut(nScanOut1743), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1744 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_16), .NorthIn(nOut27_15), .SouthIn(nOut27_17), .EastIn(nOut28_16), .WestIn(nOut26_16), .ScanIn(nScanOut1745), .ScanOut(nScanOut1744), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1745 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_17), .NorthIn(nOut27_16), .SouthIn(nOut27_18), .EastIn(nOut28_17), .WestIn(nOut26_17), .ScanIn(nScanOut1746), .ScanOut(nScanOut1745), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1746 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_18), .NorthIn(nOut27_17), .SouthIn(nOut27_19), .EastIn(nOut28_18), .WestIn(nOut26_18), .ScanIn(nScanOut1747), .ScanOut(nScanOut1746), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1747 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_19), .NorthIn(nOut27_18), .SouthIn(nOut27_20), .EastIn(nOut28_19), .WestIn(nOut26_19), .ScanIn(nScanOut1748), .ScanOut(nScanOut1747), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1748 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_20), .NorthIn(nOut27_19), .SouthIn(nOut27_21), .EastIn(nOut28_20), .WestIn(nOut26_20), .ScanIn(nScanOut1749), .ScanOut(nScanOut1748), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1749 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_21), .NorthIn(nOut27_20), .SouthIn(nOut27_22), .EastIn(nOut28_21), .WestIn(nOut26_21), .ScanIn(nScanOut1750), .ScanOut(nScanOut1749), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1750 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_22), .NorthIn(nOut27_21), .SouthIn(nOut27_23), .EastIn(nOut28_22), .WestIn(nOut26_22), .ScanIn(nScanOut1751), .ScanOut(nScanOut1750), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1751 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_23), .NorthIn(nOut27_22), .SouthIn(nOut27_24), .EastIn(nOut28_23), .WestIn(nOut26_23), .ScanIn(nScanOut1752), .ScanOut(nScanOut1751), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1752 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_24), .NorthIn(nOut27_23), .SouthIn(nOut27_25), .EastIn(nOut28_24), .WestIn(nOut26_24), .ScanIn(nScanOut1753), .ScanOut(nScanOut1752), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1753 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_25), .NorthIn(nOut27_24), .SouthIn(nOut27_26), .EastIn(nOut28_25), .WestIn(nOut26_25), .ScanIn(nScanOut1754), .ScanOut(nScanOut1753), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1754 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_26), .NorthIn(nOut27_25), .SouthIn(nOut27_27), .EastIn(nOut28_26), .WestIn(nOut26_26), .ScanIn(nScanOut1755), .ScanOut(nScanOut1754), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1755 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_27), .NorthIn(nOut27_26), .SouthIn(nOut27_28), .EastIn(nOut28_27), .WestIn(nOut26_27), .ScanIn(nScanOut1756), .ScanOut(nScanOut1755), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1756 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_28), .NorthIn(nOut27_27), .SouthIn(nOut27_29), .EastIn(nOut28_28), .WestIn(nOut26_28), .ScanIn(nScanOut1757), .ScanOut(nScanOut1756), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1757 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_29), .NorthIn(nOut27_28), .SouthIn(nOut27_30), .EastIn(nOut28_29), .WestIn(nOut26_29), .ScanIn(nScanOut1758), .ScanOut(nScanOut1757), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1758 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_30), .NorthIn(nOut27_29), .SouthIn(nOut27_31), .EastIn(nOut28_30), .WestIn(nOut26_30), .ScanIn(nScanOut1759), .ScanOut(nScanOut1758), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1759 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_31), .NorthIn(nOut27_30), .SouthIn(nOut27_32), .EastIn(nOut28_31), .WestIn(nOut26_31), .ScanIn(nScanOut1760), .ScanOut(nScanOut1759), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1760 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_32), .NorthIn(nOut27_31), .SouthIn(nOut27_33), .EastIn(nOut28_32), .WestIn(nOut26_32), .ScanIn(nScanOut1761), .ScanOut(nScanOut1760), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1761 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_33), .NorthIn(nOut27_32), .SouthIn(nOut27_34), .EastIn(nOut28_33), .WestIn(nOut26_33), .ScanIn(nScanOut1762), .ScanOut(nScanOut1761), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1762 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_34), .NorthIn(nOut27_33), .SouthIn(nOut27_35), .EastIn(nOut28_34), .WestIn(nOut26_34), .ScanIn(nScanOut1763), .ScanOut(nScanOut1762), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1763 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_35), .NorthIn(nOut27_34), .SouthIn(nOut27_36), .EastIn(nOut28_35), .WestIn(nOut26_35), .ScanIn(nScanOut1764), .ScanOut(nScanOut1763), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1764 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_36), .NorthIn(nOut27_35), .SouthIn(nOut27_37), .EastIn(nOut28_36), .WestIn(nOut26_36), .ScanIn(nScanOut1765), .ScanOut(nScanOut1764), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1765 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_37), .NorthIn(nOut27_36), .SouthIn(nOut27_38), .EastIn(nOut28_37), .WestIn(nOut26_37), .ScanIn(nScanOut1766), .ScanOut(nScanOut1765), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1766 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_38), .NorthIn(nOut27_37), .SouthIn(nOut27_39), .EastIn(nOut28_38), .WestIn(nOut26_38), .ScanIn(nScanOut1767), .ScanOut(nScanOut1766), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1767 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_39), .NorthIn(nOut27_38), .SouthIn(nOut27_40), .EastIn(nOut28_39), .WestIn(nOut26_39), .ScanIn(nScanOut1768), .ScanOut(nScanOut1767), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1768 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_40), .NorthIn(nOut27_39), .SouthIn(nOut27_41), .EastIn(nOut28_40), .WestIn(nOut26_40), .ScanIn(nScanOut1769), .ScanOut(nScanOut1768), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1769 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_41), .NorthIn(nOut27_40), .SouthIn(nOut27_42), .EastIn(nOut28_41), .WestIn(nOut26_41), .ScanIn(nScanOut1770), .ScanOut(nScanOut1769), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1770 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_42), .NorthIn(nOut27_41), .SouthIn(nOut27_43), .EastIn(nOut28_42), .WestIn(nOut26_42), .ScanIn(nScanOut1771), .ScanOut(nScanOut1770), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1771 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_43), .NorthIn(nOut27_42), .SouthIn(nOut27_44), .EastIn(nOut28_43), .WestIn(nOut26_43), .ScanIn(nScanOut1772), .ScanOut(nScanOut1771), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1772 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_44), .NorthIn(nOut27_43), .SouthIn(nOut27_45), .EastIn(nOut28_44), .WestIn(nOut26_44), .ScanIn(nScanOut1773), .ScanOut(nScanOut1772), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1773 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_45), .NorthIn(nOut27_44), .SouthIn(nOut27_46), .EastIn(nOut28_45), .WestIn(nOut26_45), .ScanIn(nScanOut1774), .ScanOut(nScanOut1773), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1774 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_46), .NorthIn(nOut27_45), .SouthIn(nOut27_47), .EastIn(nOut28_46), .WestIn(nOut26_46), .ScanIn(nScanOut1775), .ScanOut(nScanOut1774), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1775 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_47), .NorthIn(nOut27_46), .SouthIn(nOut27_48), .EastIn(nOut28_47), .WestIn(nOut26_47), .ScanIn(nScanOut1776), .ScanOut(nScanOut1775), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1776 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_48), .NorthIn(nOut27_47), .SouthIn(nOut27_49), .EastIn(nOut28_48), .WestIn(nOut26_48), .ScanIn(nScanOut1777), .ScanOut(nScanOut1776), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1777 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_49), .NorthIn(nOut27_48), .SouthIn(nOut27_50), .EastIn(nOut28_49), .WestIn(nOut26_49), .ScanIn(nScanOut1778), .ScanOut(nScanOut1777), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1778 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_50), .NorthIn(nOut27_49), .SouthIn(nOut27_51), .EastIn(nOut28_50), .WestIn(nOut26_50), .ScanIn(nScanOut1779), .ScanOut(nScanOut1778), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1779 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_51), .NorthIn(nOut27_50), .SouthIn(nOut27_52), .EastIn(nOut28_51), .WestIn(nOut26_51), .ScanIn(nScanOut1780), .ScanOut(nScanOut1779), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1780 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_52), .NorthIn(nOut27_51), .SouthIn(nOut27_53), .EastIn(nOut28_52), .WestIn(nOut26_52), .ScanIn(nScanOut1781), .ScanOut(nScanOut1780), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1781 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_53), .NorthIn(nOut27_52), .SouthIn(nOut27_54), .EastIn(nOut28_53), .WestIn(nOut26_53), .ScanIn(nScanOut1782), .ScanOut(nScanOut1781), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1782 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_54), .NorthIn(nOut27_53), .SouthIn(nOut27_55), .EastIn(nOut28_54), .WestIn(nOut26_54), .ScanIn(nScanOut1783), .ScanOut(nScanOut1782), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1783 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_55), .NorthIn(nOut27_54), .SouthIn(nOut27_56), .EastIn(nOut28_55), .WestIn(nOut26_55), .ScanIn(nScanOut1784), .ScanOut(nScanOut1783), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1784 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_56), .NorthIn(nOut27_55), .SouthIn(nOut27_57), .EastIn(nOut28_56), .WestIn(nOut26_56), .ScanIn(nScanOut1785), .ScanOut(nScanOut1784), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1785 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_57), .NorthIn(nOut27_56), .SouthIn(nOut27_58), .EastIn(nOut28_57), .WestIn(nOut26_57), .ScanIn(nScanOut1786), .ScanOut(nScanOut1785), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1786 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_58), .NorthIn(nOut27_57), .SouthIn(nOut27_59), .EastIn(nOut28_58), .WestIn(nOut26_58), .ScanIn(nScanOut1787), .ScanOut(nScanOut1786), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1787 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_59), .NorthIn(nOut27_58), .SouthIn(nOut27_60), .EastIn(nOut28_59), .WestIn(nOut26_59), .ScanIn(nScanOut1788), .ScanOut(nScanOut1787), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1788 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_60), .NorthIn(nOut27_59), .SouthIn(nOut27_61), .EastIn(nOut28_60), .WestIn(nOut26_60), .ScanIn(nScanOut1789), .ScanOut(nScanOut1788), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1789 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_61), .NorthIn(nOut27_60), .SouthIn(nOut27_62), .EastIn(nOut28_61), .WestIn(nOut26_61), .ScanIn(nScanOut1790), .ScanOut(nScanOut1789), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1790 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut27_62), .NorthIn(nOut27_61), .SouthIn(nOut27_63), .EastIn(nOut28_62), .WestIn(nOut26_62), .ScanIn(nScanOut1791), .ScanOut(nScanOut1790), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1791 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut27_63), .ScanIn(nScanOut1792), .ScanOut(nScanOut1791), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1792 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut28_0), .ScanIn(nScanOut1793), .ScanOut(nScanOut1792), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1793 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_1), .NorthIn(nOut28_0), .SouthIn(nOut28_2), .EastIn(nOut29_1), .WestIn(nOut27_1), .ScanIn(nScanOut1794), .ScanOut(nScanOut1793), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1794 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_2), .NorthIn(nOut28_1), .SouthIn(nOut28_3), .EastIn(nOut29_2), .WestIn(nOut27_2), .ScanIn(nScanOut1795), .ScanOut(nScanOut1794), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1795 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_3), .NorthIn(nOut28_2), .SouthIn(nOut28_4), .EastIn(nOut29_3), .WestIn(nOut27_3), .ScanIn(nScanOut1796), .ScanOut(nScanOut1795), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1796 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_4), .NorthIn(nOut28_3), .SouthIn(nOut28_5), .EastIn(nOut29_4), .WestIn(nOut27_4), .ScanIn(nScanOut1797), .ScanOut(nScanOut1796), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1797 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_5), .NorthIn(nOut28_4), .SouthIn(nOut28_6), .EastIn(nOut29_5), .WestIn(nOut27_5), .ScanIn(nScanOut1798), .ScanOut(nScanOut1797), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1798 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_6), .NorthIn(nOut28_5), .SouthIn(nOut28_7), .EastIn(nOut29_6), .WestIn(nOut27_6), .ScanIn(nScanOut1799), .ScanOut(nScanOut1798), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1799 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_7), .NorthIn(nOut28_6), .SouthIn(nOut28_8), .EastIn(nOut29_7), .WestIn(nOut27_7), .ScanIn(nScanOut1800), .ScanOut(nScanOut1799), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1800 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_8), .NorthIn(nOut28_7), .SouthIn(nOut28_9), .EastIn(nOut29_8), .WestIn(nOut27_8), .ScanIn(nScanOut1801), .ScanOut(nScanOut1800), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1801 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_9), .NorthIn(nOut28_8), .SouthIn(nOut28_10), .EastIn(nOut29_9), .WestIn(nOut27_9), .ScanIn(nScanOut1802), .ScanOut(nScanOut1801), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1802 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_10), .NorthIn(nOut28_9), .SouthIn(nOut28_11), .EastIn(nOut29_10), .WestIn(nOut27_10), .ScanIn(nScanOut1803), .ScanOut(nScanOut1802), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1803 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_11), .NorthIn(nOut28_10), .SouthIn(nOut28_12), .EastIn(nOut29_11), .WestIn(nOut27_11), .ScanIn(nScanOut1804), .ScanOut(nScanOut1803), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1804 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_12), .NorthIn(nOut28_11), .SouthIn(nOut28_13), .EastIn(nOut29_12), .WestIn(nOut27_12), .ScanIn(nScanOut1805), .ScanOut(nScanOut1804), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1805 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_13), .NorthIn(nOut28_12), .SouthIn(nOut28_14), .EastIn(nOut29_13), .WestIn(nOut27_13), .ScanIn(nScanOut1806), .ScanOut(nScanOut1805), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1806 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_14), .NorthIn(nOut28_13), .SouthIn(nOut28_15), .EastIn(nOut29_14), .WestIn(nOut27_14), .ScanIn(nScanOut1807), .ScanOut(nScanOut1806), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1807 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_15), .NorthIn(nOut28_14), .SouthIn(nOut28_16), .EastIn(nOut29_15), .WestIn(nOut27_15), .ScanIn(nScanOut1808), .ScanOut(nScanOut1807), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1808 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_16), .NorthIn(nOut28_15), .SouthIn(nOut28_17), .EastIn(nOut29_16), .WestIn(nOut27_16), .ScanIn(nScanOut1809), .ScanOut(nScanOut1808), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1809 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_17), .NorthIn(nOut28_16), .SouthIn(nOut28_18), .EastIn(nOut29_17), .WestIn(nOut27_17), .ScanIn(nScanOut1810), .ScanOut(nScanOut1809), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1810 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_18), .NorthIn(nOut28_17), .SouthIn(nOut28_19), .EastIn(nOut29_18), .WestIn(nOut27_18), .ScanIn(nScanOut1811), .ScanOut(nScanOut1810), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1811 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_19), .NorthIn(nOut28_18), .SouthIn(nOut28_20), .EastIn(nOut29_19), .WestIn(nOut27_19), .ScanIn(nScanOut1812), .ScanOut(nScanOut1811), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1812 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_20), .NorthIn(nOut28_19), .SouthIn(nOut28_21), .EastIn(nOut29_20), .WestIn(nOut27_20), .ScanIn(nScanOut1813), .ScanOut(nScanOut1812), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1813 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_21), .NorthIn(nOut28_20), .SouthIn(nOut28_22), .EastIn(nOut29_21), .WestIn(nOut27_21), .ScanIn(nScanOut1814), .ScanOut(nScanOut1813), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1814 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_22), .NorthIn(nOut28_21), .SouthIn(nOut28_23), .EastIn(nOut29_22), .WestIn(nOut27_22), .ScanIn(nScanOut1815), .ScanOut(nScanOut1814), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1815 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_23), .NorthIn(nOut28_22), .SouthIn(nOut28_24), .EastIn(nOut29_23), .WestIn(nOut27_23), .ScanIn(nScanOut1816), .ScanOut(nScanOut1815), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1816 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_24), .NorthIn(nOut28_23), .SouthIn(nOut28_25), .EastIn(nOut29_24), .WestIn(nOut27_24), .ScanIn(nScanOut1817), .ScanOut(nScanOut1816), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1817 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_25), .NorthIn(nOut28_24), .SouthIn(nOut28_26), .EastIn(nOut29_25), .WestIn(nOut27_25), .ScanIn(nScanOut1818), .ScanOut(nScanOut1817), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1818 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_26), .NorthIn(nOut28_25), .SouthIn(nOut28_27), .EastIn(nOut29_26), .WestIn(nOut27_26), .ScanIn(nScanOut1819), .ScanOut(nScanOut1818), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1819 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_27), .NorthIn(nOut28_26), .SouthIn(nOut28_28), .EastIn(nOut29_27), .WestIn(nOut27_27), .ScanIn(nScanOut1820), .ScanOut(nScanOut1819), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1820 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_28), .NorthIn(nOut28_27), .SouthIn(nOut28_29), .EastIn(nOut29_28), .WestIn(nOut27_28), .ScanIn(nScanOut1821), .ScanOut(nScanOut1820), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1821 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_29), .NorthIn(nOut28_28), .SouthIn(nOut28_30), .EastIn(nOut29_29), .WestIn(nOut27_29), .ScanIn(nScanOut1822), .ScanOut(nScanOut1821), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1822 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_30), .NorthIn(nOut28_29), .SouthIn(nOut28_31), .EastIn(nOut29_30), .WestIn(nOut27_30), .ScanIn(nScanOut1823), .ScanOut(nScanOut1822), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1823 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_31), .NorthIn(nOut28_30), .SouthIn(nOut28_32), .EastIn(nOut29_31), .WestIn(nOut27_31), .ScanIn(nScanOut1824), .ScanOut(nScanOut1823), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1824 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_32), .NorthIn(nOut28_31), .SouthIn(nOut28_33), .EastIn(nOut29_32), .WestIn(nOut27_32), .ScanIn(nScanOut1825), .ScanOut(nScanOut1824), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1825 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_33), .NorthIn(nOut28_32), .SouthIn(nOut28_34), .EastIn(nOut29_33), .WestIn(nOut27_33), .ScanIn(nScanOut1826), .ScanOut(nScanOut1825), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1826 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_34), .NorthIn(nOut28_33), .SouthIn(nOut28_35), .EastIn(nOut29_34), .WestIn(nOut27_34), .ScanIn(nScanOut1827), .ScanOut(nScanOut1826), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1827 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_35), .NorthIn(nOut28_34), .SouthIn(nOut28_36), .EastIn(nOut29_35), .WestIn(nOut27_35), .ScanIn(nScanOut1828), .ScanOut(nScanOut1827), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1828 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_36), .NorthIn(nOut28_35), .SouthIn(nOut28_37), .EastIn(nOut29_36), .WestIn(nOut27_36), .ScanIn(nScanOut1829), .ScanOut(nScanOut1828), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1829 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_37), .NorthIn(nOut28_36), .SouthIn(nOut28_38), .EastIn(nOut29_37), .WestIn(nOut27_37), .ScanIn(nScanOut1830), .ScanOut(nScanOut1829), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1830 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_38), .NorthIn(nOut28_37), .SouthIn(nOut28_39), .EastIn(nOut29_38), .WestIn(nOut27_38), .ScanIn(nScanOut1831), .ScanOut(nScanOut1830), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1831 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_39), .NorthIn(nOut28_38), .SouthIn(nOut28_40), .EastIn(nOut29_39), .WestIn(nOut27_39), .ScanIn(nScanOut1832), .ScanOut(nScanOut1831), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1832 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_40), .NorthIn(nOut28_39), .SouthIn(nOut28_41), .EastIn(nOut29_40), .WestIn(nOut27_40), .ScanIn(nScanOut1833), .ScanOut(nScanOut1832), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1833 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_41), .NorthIn(nOut28_40), .SouthIn(nOut28_42), .EastIn(nOut29_41), .WestIn(nOut27_41), .ScanIn(nScanOut1834), .ScanOut(nScanOut1833), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1834 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_42), .NorthIn(nOut28_41), .SouthIn(nOut28_43), .EastIn(nOut29_42), .WestIn(nOut27_42), .ScanIn(nScanOut1835), .ScanOut(nScanOut1834), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1835 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_43), .NorthIn(nOut28_42), .SouthIn(nOut28_44), .EastIn(nOut29_43), .WestIn(nOut27_43), .ScanIn(nScanOut1836), .ScanOut(nScanOut1835), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1836 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_44), .NorthIn(nOut28_43), .SouthIn(nOut28_45), .EastIn(nOut29_44), .WestIn(nOut27_44), .ScanIn(nScanOut1837), .ScanOut(nScanOut1836), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1837 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_45), .NorthIn(nOut28_44), .SouthIn(nOut28_46), .EastIn(nOut29_45), .WestIn(nOut27_45), .ScanIn(nScanOut1838), .ScanOut(nScanOut1837), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1838 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_46), .NorthIn(nOut28_45), .SouthIn(nOut28_47), .EastIn(nOut29_46), .WestIn(nOut27_46), .ScanIn(nScanOut1839), .ScanOut(nScanOut1838), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1839 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_47), .NorthIn(nOut28_46), .SouthIn(nOut28_48), .EastIn(nOut29_47), .WestIn(nOut27_47), .ScanIn(nScanOut1840), .ScanOut(nScanOut1839), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1840 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_48), .NorthIn(nOut28_47), .SouthIn(nOut28_49), .EastIn(nOut29_48), .WestIn(nOut27_48), .ScanIn(nScanOut1841), .ScanOut(nScanOut1840), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1841 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_49), .NorthIn(nOut28_48), .SouthIn(nOut28_50), .EastIn(nOut29_49), .WestIn(nOut27_49), .ScanIn(nScanOut1842), .ScanOut(nScanOut1841), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1842 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_50), .NorthIn(nOut28_49), .SouthIn(nOut28_51), .EastIn(nOut29_50), .WestIn(nOut27_50), .ScanIn(nScanOut1843), .ScanOut(nScanOut1842), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1843 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_51), .NorthIn(nOut28_50), .SouthIn(nOut28_52), .EastIn(nOut29_51), .WestIn(nOut27_51), .ScanIn(nScanOut1844), .ScanOut(nScanOut1843), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1844 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_52), .NorthIn(nOut28_51), .SouthIn(nOut28_53), .EastIn(nOut29_52), .WestIn(nOut27_52), .ScanIn(nScanOut1845), .ScanOut(nScanOut1844), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1845 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_53), .NorthIn(nOut28_52), .SouthIn(nOut28_54), .EastIn(nOut29_53), .WestIn(nOut27_53), .ScanIn(nScanOut1846), .ScanOut(nScanOut1845), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1846 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_54), .NorthIn(nOut28_53), .SouthIn(nOut28_55), .EastIn(nOut29_54), .WestIn(nOut27_54), .ScanIn(nScanOut1847), .ScanOut(nScanOut1846), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1847 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_55), .NorthIn(nOut28_54), .SouthIn(nOut28_56), .EastIn(nOut29_55), .WestIn(nOut27_55), .ScanIn(nScanOut1848), .ScanOut(nScanOut1847), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1848 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_56), .NorthIn(nOut28_55), .SouthIn(nOut28_57), .EastIn(nOut29_56), .WestIn(nOut27_56), .ScanIn(nScanOut1849), .ScanOut(nScanOut1848), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1849 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_57), .NorthIn(nOut28_56), .SouthIn(nOut28_58), .EastIn(nOut29_57), .WestIn(nOut27_57), .ScanIn(nScanOut1850), .ScanOut(nScanOut1849), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1850 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_58), .NorthIn(nOut28_57), .SouthIn(nOut28_59), .EastIn(nOut29_58), .WestIn(nOut27_58), .ScanIn(nScanOut1851), .ScanOut(nScanOut1850), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1851 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_59), .NorthIn(nOut28_58), .SouthIn(nOut28_60), .EastIn(nOut29_59), .WestIn(nOut27_59), .ScanIn(nScanOut1852), .ScanOut(nScanOut1851), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1852 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_60), .NorthIn(nOut28_59), .SouthIn(nOut28_61), .EastIn(nOut29_60), .WestIn(nOut27_60), .ScanIn(nScanOut1853), .ScanOut(nScanOut1852), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1853 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_61), .NorthIn(nOut28_60), .SouthIn(nOut28_62), .EastIn(nOut29_61), .WestIn(nOut27_61), .ScanIn(nScanOut1854), .ScanOut(nScanOut1853), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1854 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut28_62), .NorthIn(nOut28_61), .SouthIn(nOut28_63), .EastIn(nOut29_62), .WestIn(nOut27_62), .ScanIn(nScanOut1855), .ScanOut(nScanOut1854), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1855 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut28_63), .ScanIn(nScanOut1856), .ScanOut(nScanOut1855), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1856 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut29_0), .ScanIn(nScanOut1857), .ScanOut(nScanOut1856), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1857 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_1), .NorthIn(nOut29_0), .SouthIn(nOut29_2), .EastIn(nOut30_1), .WestIn(nOut28_1), .ScanIn(nScanOut1858), .ScanOut(nScanOut1857), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1858 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_2), .NorthIn(nOut29_1), .SouthIn(nOut29_3), .EastIn(nOut30_2), .WestIn(nOut28_2), .ScanIn(nScanOut1859), .ScanOut(nScanOut1858), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1859 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_3), .NorthIn(nOut29_2), .SouthIn(nOut29_4), .EastIn(nOut30_3), .WestIn(nOut28_3), .ScanIn(nScanOut1860), .ScanOut(nScanOut1859), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1860 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_4), .NorthIn(nOut29_3), .SouthIn(nOut29_5), .EastIn(nOut30_4), .WestIn(nOut28_4), .ScanIn(nScanOut1861), .ScanOut(nScanOut1860), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1861 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_5), .NorthIn(nOut29_4), .SouthIn(nOut29_6), .EastIn(nOut30_5), .WestIn(nOut28_5), .ScanIn(nScanOut1862), .ScanOut(nScanOut1861), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1862 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_6), .NorthIn(nOut29_5), .SouthIn(nOut29_7), .EastIn(nOut30_6), .WestIn(nOut28_6), .ScanIn(nScanOut1863), .ScanOut(nScanOut1862), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1863 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_7), .NorthIn(nOut29_6), .SouthIn(nOut29_8), .EastIn(nOut30_7), .WestIn(nOut28_7), .ScanIn(nScanOut1864), .ScanOut(nScanOut1863), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1864 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_8), .NorthIn(nOut29_7), .SouthIn(nOut29_9), .EastIn(nOut30_8), .WestIn(nOut28_8), .ScanIn(nScanOut1865), .ScanOut(nScanOut1864), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1865 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_9), .NorthIn(nOut29_8), .SouthIn(nOut29_10), .EastIn(nOut30_9), .WestIn(nOut28_9), .ScanIn(nScanOut1866), .ScanOut(nScanOut1865), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1866 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_10), .NorthIn(nOut29_9), .SouthIn(nOut29_11), .EastIn(nOut30_10), .WestIn(nOut28_10), .ScanIn(nScanOut1867), .ScanOut(nScanOut1866), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1867 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_11), .NorthIn(nOut29_10), .SouthIn(nOut29_12), .EastIn(nOut30_11), .WestIn(nOut28_11), .ScanIn(nScanOut1868), .ScanOut(nScanOut1867), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1868 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_12), .NorthIn(nOut29_11), .SouthIn(nOut29_13), .EastIn(nOut30_12), .WestIn(nOut28_12), .ScanIn(nScanOut1869), .ScanOut(nScanOut1868), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1869 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_13), .NorthIn(nOut29_12), .SouthIn(nOut29_14), .EastIn(nOut30_13), .WestIn(nOut28_13), .ScanIn(nScanOut1870), .ScanOut(nScanOut1869), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1870 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_14), .NorthIn(nOut29_13), .SouthIn(nOut29_15), .EastIn(nOut30_14), .WestIn(nOut28_14), .ScanIn(nScanOut1871), .ScanOut(nScanOut1870), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1871 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_15), .NorthIn(nOut29_14), .SouthIn(nOut29_16), .EastIn(nOut30_15), .WestIn(nOut28_15), .ScanIn(nScanOut1872), .ScanOut(nScanOut1871), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1872 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_16), .NorthIn(nOut29_15), .SouthIn(nOut29_17), .EastIn(nOut30_16), .WestIn(nOut28_16), .ScanIn(nScanOut1873), .ScanOut(nScanOut1872), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1873 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_17), .NorthIn(nOut29_16), .SouthIn(nOut29_18), .EastIn(nOut30_17), .WestIn(nOut28_17), .ScanIn(nScanOut1874), .ScanOut(nScanOut1873), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1874 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_18), .NorthIn(nOut29_17), .SouthIn(nOut29_19), .EastIn(nOut30_18), .WestIn(nOut28_18), .ScanIn(nScanOut1875), .ScanOut(nScanOut1874), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1875 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_19), .NorthIn(nOut29_18), .SouthIn(nOut29_20), .EastIn(nOut30_19), .WestIn(nOut28_19), .ScanIn(nScanOut1876), .ScanOut(nScanOut1875), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1876 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_20), .NorthIn(nOut29_19), .SouthIn(nOut29_21), .EastIn(nOut30_20), .WestIn(nOut28_20), .ScanIn(nScanOut1877), .ScanOut(nScanOut1876), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1877 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_21), .NorthIn(nOut29_20), .SouthIn(nOut29_22), .EastIn(nOut30_21), .WestIn(nOut28_21), .ScanIn(nScanOut1878), .ScanOut(nScanOut1877), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1878 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_22), .NorthIn(nOut29_21), .SouthIn(nOut29_23), .EastIn(nOut30_22), .WestIn(nOut28_22), .ScanIn(nScanOut1879), .ScanOut(nScanOut1878), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1879 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_23), .NorthIn(nOut29_22), .SouthIn(nOut29_24), .EastIn(nOut30_23), .WestIn(nOut28_23), .ScanIn(nScanOut1880), .ScanOut(nScanOut1879), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1880 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_24), .NorthIn(nOut29_23), .SouthIn(nOut29_25), .EastIn(nOut30_24), .WestIn(nOut28_24), .ScanIn(nScanOut1881), .ScanOut(nScanOut1880), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1881 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_25), .NorthIn(nOut29_24), .SouthIn(nOut29_26), .EastIn(nOut30_25), .WestIn(nOut28_25), .ScanIn(nScanOut1882), .ScanOut(nScanOut1881), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1882 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_26), .NorthIn(nOut29_25), .SouthIn(nOut29_27), .EastIn(nOut30_26), .WestIn(nOut28_26), .ScanIn(nScanOut1883), .ScanOut(nScanOut1882), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1883 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_27), .NorthIn(nOut29_26), .SouthIn(nOut29_28), .EastIn(nOut30_27), .WestIn(nOut28_27), .ScanIn(nScanOut1884), .ScanOut(nScanOut1883), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1884 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_28), .NorthIn(nOut29_27), .SouthIn(nOut29_29), .EastIn(nOut30_28), .WestIn(nOut28_28), .ScanIn(nScanOut1885), .ScanOut(nScanOut1884), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1885 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_29), .NorthIn(nOut29_28), .SouthIn(nOut29_30), .EastIn(nOut30_29), .WestIn(nOut28_29), .ScanIn(nScanOut1886), .ScanOut(nScanOut1885), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1886 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_30), .NorthIn(nOut29_29), .SouthIn(nOut29_31), .EastIn(nOut30_30), .WestIn(nOut28_30), .ScanIn(nScanOut1887), .ScanOut(nScanOut1886), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1887 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_31), .NorthIn(nOut29_30), .SouthIn(nOut29_32), .EastIn(nOut30_31), .WestIn(nOut28_31), .ScanIn(nScanOut1888), .ScanOut(nScanOut1887), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1888 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_32), .NorthIn(nOut29_31), .SouthIn(nOut29_33), .EastIn(nOut30_32), .WestIn(nOut28_32), .ScanIn(nScanOut1889), .ScanOut(nScanOut1888), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1889 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_33), .NorthIn(nOut29_32), .SouthIn(nOut29_34), .EastIn(nOut30_33), .WestIn(nOut28_33), .ScanIn(nScanOut1890), .ScanOut(nScanOut1889), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1890 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_34), .NorthIn(nOut29_33), .SouthIn(nOut29_35), .EastIn(nOut30_34), .WestIn(nOut28_34), .ScanIn(nScanOut1891), .ScanOut(nScanOut1890), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1891 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_35), .NorthIn(nOut29_34), .SouthIn(nOut29_36), .EastIn(nOut30_35), .WestIn(nOut28_35), .ScanIn(nScanOut1892), .ScanOut(nScanOut1891), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1892 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_36), .NorthIn(nOut29_35), .SouthIn(nOut29_37), .EastIn(nOut30_36), .WestIn(nOut28_36), .ScanIn(nScanOut1893), .ScanOut(nScanOut1892), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1893 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_37), .NorthIn(nOut29_36), .SouthIn(nOut29_38), .EastIn(nOut30_37), .WestIn(nOut28_37), .ScanIn(nScanOut1894), .ScanOut(nScanOut1893), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1894 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_38), .NorthIn(nOut29_37), .SouthIn(nOut29_39), .EastIn(nOut30_38), .WestIn(nOut28_38), .ScanIn(nScanOut1895), .ScanOut(nScanOut1894), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1895 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_39), .NorthIn(nOut29_38), .SouthIn(nOut29_40), .EastIn(nOut30_39), .WestIn(nOut28_39), .ScanIn(nScanOut1896), .ScanOut(nScanOut1895), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1896 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_40), .NorthIn(nOut29_39), .SouthIn(nOut29_41), .EastIn(nOut30_40), .WestIn(nOut28_40), .ScanIn(nScanOut1897), .ScanOut(nScanOut1896), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1897 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_41), .NorthIn(nOut29_40), .SouthIn(nOut29_42), .EastIn(nOut30_41), .WestIn(nOut28_41), .ScanIn(nScanOut1898), .ScanOut(nScanOut1897), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1898 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_42), .NorthIn(nOut29_41), .SouthIn(nOut29_43), .EastIn(nOut30_42), .WestIn(nOut28_42), .ScanIn(nScanOut1899), .ScanOut(nScanOut1898), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1899 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_43), .NorthIn(nOut29_42), .SouthIn(nOut29_44), .EastIn(nOut30_43), .WestIn(nOut28_43), .ScanIn(nScanOut1900), .ScanOut(nScanOut1899), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1900 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_44), .NorthIn(nOut29_43), .SouthIn(nOut29_45), .EastIn(nOut30_44), .WestIn(nOut28_44), .ScanIn(nScanOut1901), .ScanOut(nScanOut1900), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1901 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_45), .NorthIn(nOut29_44), .SouthIn(nOut29_46), .EastIn(nOut30_45), .WestIn(nOut28_45), .ScanIn(nScanOut1902), .ScanOut(nScanOut1901), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1902 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_46), .NorthIn(nOut29_45), .SouthIn(nOut29_47), .EastIn(nOut30_46), .WestIn(nOut28_46), .ScanIn(nScanOut1903), .ScanOut(nScanOut1902), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1903 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_47), .NorthIn(nOut29_46), .SouthIn(nOut29_48), .EastIn(nOut30_47), .WestIn(nOut28_47), .ScanIn(nScanOut1904), .ScanOut(nScanOut1903), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1904 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_48), .NorthIn(nOut29_47), .SouthIn(nOut29_49), .EastIn(nOut30_48), .WestIn(nOut28_48), .ScanIn(nScanOut1905), .ScanOut(nScanOut1904), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1905 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_49), .NorthIn(nOut29_48), .SouthIn(nOut29_50), .EastIn(nOut30_49), .WestIn(nOut28_49), .ScanIn(nScanOut1906), .ScanOut(nScanOut1905), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1906 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_50), .NorthIn(nOut29_49), .SouthIn(nOut29_51), .EastIn(nOut30_50), .WestIn(nOut28_50), .ScanIn(nScanOut1907), .ScanOut(nScanOut1906), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1907 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_51), .NorthIn(nOut29_50), .SouthIn(nOut29_52), .EastIn(nOut30_51), .WestIn(nOut28_51), .ScanIn(nScanOut1908), .ScanOut(nScanOut1907), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1908 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_52), .NorthIn(nOut29_51), .SouthIn(nOut29_53), .EastIn(nOut30_52), .WestIn(nOut28_52), .ScanIn(nScanOut1909), .ScanOut(nScanOut1908), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1909 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_53), .NorthIn(nOut29_52), .SouthIn(nOut29_54), .EastIn(nOut30_53), .WestIn(nOut28_53), .ScanIn(nScanOut1910), .ScanOut(nScanOut1909), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1910 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_54), .NorthIn(nOut29_53), .SouthIn(nOut29_55), .EastIn(nOut30_54), .WestIn(nOut28_54), .ScanIn(nScanOut1911), .ScanOut(nScanOut1910), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1911 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_55), .NorthIn(nOut29_54), .SouthIn(nOut29_56), .EastIn(nOut30_55), .WestIn(nOut28_55), .ScanIn(nScanOut1912), .ScanOut(nScanOut1911), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1912 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_56), .NorthIn(nOut29_55), .SouthIn(nOut29_57), .EastIn(nOut30_56), .WestIn(nOut28_56), .ScanIn(nScanOut1913), .ScanOut(nScanOut1912), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1913 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_57), .NorthIn(nOut29_56), .SouthIn(nOut29_58), .EastIn(nOut30_57), .WestIn(nOut28_57), .ScanIn(nScanOut1914), .ScanOut(nScanOut1913), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1914 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_58), .NorthIn(nOut29_57), .SouthIn(nOut29_59), .EastIn(nOut30_58), .WestIn(nOut28_58), .ScanIn(nScanOut1915), .ScanOut(nScanOut1914), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1915 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_59), .NorthIn(nOut29_58), .SouthIn(nOut29_60), .EastIn(nOut30_59), .WestIn(nOut28_59), .ScanIn(nScanOut1916), .ScanOut(nScanOut1915), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1916 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_60), .NorthIn(nOut29_59), .SouthIn(nOut29_61), .EastIn(nOut30_60), .WestIn(nOut28_60), .ScanIn(nScanOut1917), .ScanOut(nScanOut1916), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1917 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_61), .NorthIn(nOut29_60), .SouthIn(nOut29_62), .EastIn(nOut30_61), .WestIn(nOut28_61), .ScanIn(nScanOut1918), .ScanOut(nScanOut1917), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1918 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut29_62), .NorthIn(nOut29_61), .SouthIn(nOut29_63), .EastIn(nOut30_62), .WestIn(nOut28_62), .ScanIn(nScanOut1919), .ScanOut(nScanOut1918), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1919 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut29_63), .ScanIn(nScanOut1920), .ScanOut(nScanOut1919), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1920 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut30_0), .ScanIn(nScanOut1921), .ScanOut(nScanOut1920), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1921 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_1), .NorthIn(nOut30_0), .SouthIn(nOut30_2), .EastIn(nOut31_1), .WestIn(nOut29_1), .ScanIn(nScanOut1922), .ScanOut(nScanOut1921), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1922 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_2), .NorthIn(nOut30_1), .SouthIn(nOut30_3), .EastIn(nOut31_2), .WestIn(nOut29_2), .ScanIn(nScanOut1923), .ScanOut(nScanOut1922), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1923 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_3), .NorthIn(nOut30_2), .SouthIn(nOut30_4), .EastIn(nOut31_3), .WestIn(nOut29_3), .ScanIn(nScanOut1924), .ScanOut(nScanOut1923), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1924 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_4), .NorthIn(nOut30_3), .SouthIn(nOut30_5), .EastIn(nOut31_4), .WestIn(nOut29_4), .ScanIn(nScanOut1925), .ScanOut(nScanOut1924), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1925 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_5), .NorthIn(nOut30_4), .SouthIn(nOut30_6), .EastIn(nOut31_5), .WestIn(nOut29_5), .ScanIn(nScanOut1926), .ScanOut(nScanOut1925), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1926 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_6), .NorthIn(nOut30_5), .SouthIn(nOut30_7), .EastIn(nOut31_6), .WestIn(nOut29_6), .ScanIn(nScanOut1927), .ScanOut(nScanOut1926), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1927 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_7), .NorthIn(nOut30_6), .SouthIn(nOut30_8), .EastIn(nOut31_7), .WestIn(nOut29_7), .ScanIn(nScanOut1928), .ScanOut(nScanOut1927), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1928 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_8), .NorthIn(nOut30_7), .SouthIn(nOut30_9), .EastIn(nOut31_8), .WestIn(nOut29_8), .ScanIn(nScanOut1929), .ScanOut(nScanOut1928), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1929 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_9), .NorthIn(nOut30_8), .SouthIn(nOut30_10), .EastIn(nOut31_9), .WestIn(nOut29_9), .ScanIn(nScanOut1930), .ScanOut(nScanOut1929), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1930 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_10), .NorthIn(nOut30_9), .SouthIn(nOut30_11), .EastIn(nOut31_10), .WestIn(nOut29_10), .ScanIn(nScanOut1931), .ScanOut(nScanOut1930), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1931 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_11), .NorthIn(nOut30_10), .SouthIn(nOut30_12), .EastIn(nOut31_11), .WestIn(nOut29_11), .ScanIn(nScanOut1932), .ScanOut(nScanOut1931), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1932 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_12), .NorthIn(nOut30_11), .SouthIn(nOut30_13), .EastIn(nOut31_12), .WestIn(nOut29_12), .ScanIn(nScanOut1933), .ScanOut(nScanOut1932), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1933 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_13), .NorthIn(nOut30_12), .SouthIn(nOut30_14), .EastIn(nOut31_13), .WestIn(nOut29_13), .ScanIn(nScanOut1934), .ScanOut(nScanOut1933), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1934 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_14), .NorthIn(nOut30_13), .SouthIn(nOut30_15), .EastIn(nOut31_14), .WestIn(nOut29_14), .ScanIn(nScanOut1935), .ScanOut(nScanOut1934), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1935 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_15), .NorthIn(nOut30_14), .SouthIn(nOut30_16), .EastIn(nOut31_15), .WestIn(nOut29_15), .ScanIn(nScanOut1936), .ScanOut(nScanOut1935), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1936 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_16), .NorthIn(nOut30_15), .SouthIn(nOut30_17), .EastIn(nOut31_16), .WestIn(nOut29_16), .ScanIn(nScanOut1937), .ScanOut(nScanOut1936), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1937 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_17), .NorthIn(nOut30_16), .SouthIn(nOut30_18), .EastIn(nOut31_17), .WestIn(nOut29_17), .ScanIn(nScanOut1938), .ScanOut(nScanOut1937), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1938 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_18), .NorthIn(nOut30_17), .SouthIn(nOut30_19), .EastIn(nOut31_18), .WestIn(nOut29_18), .ScanIn(nScanOut1939), .ScanOut(nScanOut1938), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1939 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_19), .NorthIn(nOut30_18), .SouthIn(nOut30_20), .EastIn(nOut31_19), .WestIn(nOut29_19), .ScanIn(nScanOut1940), .ScanOut(nScanOut1939), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1940 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_20), .NorthIn(nOut30_19), .SouthIn(nOut30_21), .EastIn(nOut31_20), .WestIn(nOut29_20), .ScanIn(nScanOut1941), .ScanOut(nScanOut1940), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1941 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_21), .NorthIn(nOut30_20), .SouthIn(nOut30_22), .EastIn(nOut31_21), .WestIn(nOut29_21), .ScanIn(nScanOut1942), .ScanOut(nScanOut1941), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1942 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_22), .NorthIn(nOut30_21), .SouthIn(nOut30_23), .EastIn(nOut31_22), .WestIn(nOut29_22), .ScanIn(nScanOut1943), .ScanOut(nScanOut1942), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1943 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_23), .NorthIn(nOut30_22), .SouthIn(nOut30_24), .EastIn(nOut31_23), .WestIn(nOut29_23), .ScanIn(nScanOut1944), .ScanOut(nScanOut1943), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1944 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_24), .NorthIn(nOut30_23), .SouthIn(nOut30_25), .EastIn(nOut31_24), .WestIn(nOut29_24), .ScanIn(nScanOut1945), .ScanOut(nScanOut1944), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1945 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_25), .NorthIn(nOut30_24), .SouthIn(nOut30_26), .EastIn(nOut31_25), .WestIn(nOut29_25), .ScanIn(nScanOut1946), .ScanOut(nScanOut1945), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1946 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_26), .NorthIn(nOut30_25), .SouthIn(nOut30_27), .EastIn(nOut31_26), .WestIn(nOut29_26), .ScanIn(nScanOut1947), .ScanOut(nScanOut1946), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1947 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_27), .NorthIn(nOut30_26), .SouthIn(nOut30_28), .EastIn(nOut31_27), .WestIn(nOut29_27), .ScanIn(nScanOut1948), .ScanOut(nScanOut1947), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1948 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_28), .NorthIn(nOut30_27), .SouthIn(nOut30_29), .EastIn(nOut31_28), .WestIn(nOut29_28), .ScanIn(nScanOut1949), .ScanOut(nScanOut1948), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1949 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_29), .NorthIn(nOut30_28), .SouthIn(nOut30_30), .EastIn(nOut31_29), .WestIn(nOut29_29), .ScanIn(nScanOut1950), .ScanOut(nScanOut1949), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1950 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_30), .NorthIn(nOut30_29), .SouthIn(nOut30_31), .EastIn(nOut31_30), .WestIn(nOut29_30), .ScanIn(nScanOut1951), .ScanOut(nScanOut1950), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1951 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_31), .NorthIn(nOut30_30), .SouthIn(nOut30_32), .EastIn(nOut31_31), .WestIn(nOut29_31), .ScanIn(nScanOut1952), .ScanOut(nScanOut1951), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1952 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_32), .NorthIn(nOut30_31), .SouthIn(nOut30_33), .EastIn(nOut31_32), .WestIn(nOut29_32), .ScanIn(nScanOut1953), .ScanOut(nScanOut1952), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1953 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_33), .NorthIn(nOut30_32), .SouthIn(nOut30_34), .EastIn(nOut31_33), .WestIn(nOut29_33), .ScanIn(nScanOut1954), .ScanOut(nScanOut1953), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1954 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_34), .NorthIn(nOut30_33), .SouthIn(nOut30_35), .EastIn(nOut31_34), .WestIn(nOut29_34), .ScanIn(nScanOut1955), .ScanOut(nScanOut1954), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1955 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_35), .NorthIn(nOut30_34), .SouthIn(nOut30_36), .EastIn(nOut31_35), .WestIn(nOut29_35), .ScanIn(nScanOut1956), .ScanOut(nScanOut1955), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1956 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_36), .NorthIn(nOut30_35), .SouthIn(nOut30_37), .EastIn(nOut31_36), .WestIn(nOut29_36), .ScanIn(nScanOut1957), .ScanOut(nScanOut1956), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1957 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_37), .NorthIn(nOut30_36), .SouthIn(nOut30_38), .EastIn(nOut31_37), .WestIn(nOut29_37), .ScanIn(nScanOut1958), .ScanOut(nScanOut1957), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1958 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_38), .NorthIn(nOut30_37), .SouthIn(nOut30_39), .EastIn(nOut31_38), .WestIn(nOut29_38), .ScanIn(nScanOut1959), .ScanOut(nScanOut1958), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1959 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_39), .NorthIn(nOut30_38), .SouthIn(nOut30_40), .EastIn(nOut31_39), .WestIn(nOut29_39), .ScanIn(nScanOut1960), .ScanOut(nScanOut1959), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1960 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_40), .NorthIn(nOut30_39), .SouthIn(nOut30_41), .EastIn(nOut31_40), .WestIn(nOut29_40), .ScanIn(nScanOut1961), .ScanOut(nScanOut1960), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1961 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_41), .NorthIn(nOut30_40), .SouthIn(nOut30_42), .EastIn(nOut31_41), .WestIn(nOut29_41), .ScanIn(nScanOut1962), .ScanOut(nScanOut1961), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1962 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_42), .NorthIn(nOut30_41), .SouthIn(nOut30_43), .EastIn(nOut31_42), .WestIn(nOut29_42), .ScanIn(nScanOut1963), .ScanOut(nScanOut1962), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1963 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_43), .NorthIn(nOut30_42), .SouthIn(nOut30_44), .EastIn(nOut31_43), .WestIn(nOut29_43), .ScanIn(nScanOut1964), .ScanOut(nScanOut1963), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1964 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_44), .NorthIn(nOut30_43), .SouthIn(nOut30_45), .EastIn(nOut31_44), .WestIn(nOut29_44), .ScanIn(nScanOut1965), .ScanOut(nScanOut1964), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1965 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_45), .NorthIn(nOut30_44), .SouthIn(nOut30_46), .EastIn(nOut31_45), .WestIn(nOut29_45), .ScanIn(nScanOut1966), .ScanOut(nScanOut1965), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1966 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_46), .NorthIn(nOut30_45), .SouthIn(nOut30_47), .EastIn(nOut31_46), .WestIn(nOut29_46), .ScanIn(nScanOut1967), .ScanOut(nScanOut1966), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1967 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_47), .NorthIn(nOut30_46), .SouthIn(nOut30_48), .EastIn(nOut31_47), .WestIn(nOut29_47), .ScanIn(nScanOut1968), .ScanOut(nScanOut1967), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1968 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_48), .NorthIn(nOut30_47), .SouthIn(nOut30_49), .EastIn(nOut31_48), .WestIn(nOut29_48), .ScanIn(nScanOut1969), .ScanOut(nScanOut1968), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1969 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_49), .NorthIn(nOut30_48), .SouthIn(nOut30_50), .EastIn(nOut31_49), .WestIn(nOut29_49), .ScanIn(nScanOut1970), .ScanOut(nScanOut1969), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1970 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_50), .NorthIn(nOut30_49), .SouthIn(nOut30_51), .EastIn(nOut31_50), .WestIn(nOut29_50), .ScanIn(nScanOut1971), .ScanOut(nScanOut1970), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1971 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_51), .NorthIn(nOut30_50), .SouthIn(nOut30_52), .EastIn(nOut31_51), .WestIn(nOut29_51), .ScanIn(nScanOut1972), .ScanOut(nScanOut1971), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1972 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_52), .NorthIn(nOut30_51), .SouthIn(nOut30_53), .EastIn(nOut31_52), .WestIn(nOut29_52), .ScanIn(nScanOut1973), .ScanOut(nScanOut1972), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1973 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_53), .NorthIn(nOut30_52), .SouthIn(nOut30_54), .EastIn(nOut31_53), .WestIn(nOut29_53), .ScanIn(nScanOut1974), .ScanOut(nScanOut1973), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1974 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_54), .NorthIn(nOut30_53), .SouthIn(nOut30_55), .EastIn(nOut31_54), .WestIn(nOut29_54), .ScanIn(nScanOut1975), .ScanOut(nScanOut1974), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1975 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_55), .NorthIn(nOut30_54), .SouthIn(nOut30_56), .EastIn(nOut31_55), .WestIn(nOut29_55), .ScanIn(nScanOut1976), .ScanOut(nScanOut1975), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1976 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_56), .NorthIn(nOut30_55), .SouthIn(nOut30_57), .EastIn(nOut31_56), .WestIn(nOut29_56), .ScanIn(nScanOut1977), .ScanOut(nScanOut1976), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1977 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_57), .NorthIn(nOut30_56), .SouthIn(nOut30_58), .EastIn(nOut31_57), .WestIn(nOut29_57), .ScanIn(nScanOut1978), .ScanOut(nScanOut1977), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1978 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_58), .NorthIn(nOut30_57), .SouthIn(nOut30_59), .EastIn(nOut31_58), .WestIn(nOut29_58), .ScanIn(nScanOut1979), .ScanOut(nScanOut1978), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1979 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_59), .NorthIn(nOut30_58), .SouthIn(nOut30_60), .EastIn(nOut31_59), .WestIn(nOut29_59), .ScanIn(nScanOut1980), .ScanOut(nScanOut1979), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1980 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_60), .NorthIn(nOut30_59), .SouthIn(nOut30_61), .EastIn(nOut31_60), .WestIn(nOut29_60), .ScanIn(nScanOut1981), .ScanOut(nScanOut1980), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1981 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_61), .NorthIn(nOut30_60), .SouthIn(nOut30_62), .EastIn(nOut31_61), .WestIn(nOut29_61), .ScanIn(nScanOut1982), .ScanOut(nScanOut1981), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_1982 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut30_62), .NorthIn(nOut30_61), .SouthIn(nOut30_63), .EastIn(nOut31_62), .WestIn(nOut29_62), .ScanIn(nScanOut1983), .ScanOut(nScanOut1982), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1983 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut30_63), .ScanIn(nScanOut1984), .ScanOut(nScanOut1983), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1984 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_0), .ScanIn(nScanOut1985), .ScanOut(nScanOut1984), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1985 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_1), .ScanIn(nScanOut1986), .ScanOut(nScanOut1985), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1986 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_2), .ScanIn(nScanOut1987), .ScanOut(nScanOut1986), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1987 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_3), .ScanIn(nScanOut1988), .ScanOut(nScanOut1987), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1988 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_4), .ScanIn(nScanOut1989), .ScanOut(nScanOut1988), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1989 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_5), .ScanIn(nScanOut1990), .ScanOut(nScanOut1989), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1990 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_6), .ScanIn(nScanOut1991), .ScanOut(nScanOut1990), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1991 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_7), .ScanIn(nScanOut1992), .ScanOut(nScanOut1991), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1992 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_8), .ScanIn(nScanOut1993), .ScanOut(nScanOut1992), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1993 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_9), .ScanIn(nScanOut1994), .ScanOut(nScanOut1993), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1994 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_10), .ScanIn(nScanOut1995), .ScanOut(nScanOut1994), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1995 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_11), .ScanIn(nScanOut1996), .ScanOut(nScanOut1995), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1996 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_12), .ScanIn(nScanOut1997), .ScanOut(nScanOut1996), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1997 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_13), .ScanIn(nScanOut1998), .ScanOut(nScanOut1997), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1998 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_14), .ScanIn(nScanOut1999), .ScanOut(nScanOut1998), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1999 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_15), .ScanIn(nScanOut2000), .ScanOut(nScanOut1999), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2000 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_16), .ScanIn(nScanOut2001), .ScanOut(nScanOut2000), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2001 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_17), .ScanIn(nScanOut2002), .ScanOut(nScanOut2001), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2002 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_18), .ScanIn(nScanOut2003), .ScanOut(nScanOut2002), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2003 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_19), .ScanIn(nScanOut2004), .ScanOut(nScanOut2003), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2004 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_20), .ScanIn(nScanOut2005), .ScanOut(nScanOut2004), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2005 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_21), .ScanIn(nScanOut2006), .ScanOut(nScanOut2005), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2006 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_22), .ScanIn(nScanOut2007), .ScanOut(nScanOut2006), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2007 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_23), .ScanIn(nScanOut2008), .ScanOut(nScanOut2007), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2008 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_24), .ScanIn(nScanOut2009), .ScanOut(nScanOut2008), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2009 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_25), .ScanIn(nScanOut2010), .ScanOut(nScanOut2009), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2010 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_26), .ScanIn(nScanOut2011), .ScanOut(nScanOut2010), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2011 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_27), .ScanIn(nScanOut2012), .ScanOut(nScanOut2011), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2012 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_28), .ScanIn(nScanOut2013), .ScanOut(nScanOut2012), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2013 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_29), .ScanIn(nScanOut2014), .ScanOut(nScanOut2013), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2014 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_30), .ScanIn(nScanOut2015), .ScanOut(nScanOut2014), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2015 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_31), .ScanIn(nScanOut2016), .ScanOut(nScanOut2015), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2016 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_32), .ScanIn(nScanOut2017), .ScanOut(nScanOut2016), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2017 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_33), .ScanIn(nScanOut2018), .ScanOut(nScanOut2017), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2018 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_34), .ScanIn(nScanOut2019), .ScanOut(nScanOut2018), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2019 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_35), .ScanIn(nScanOut2020), .ScanOut(nScanOut2019), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2020 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_36), .ScanIn(nScanOut2021), .ScanOut(nScanOut2020), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2021 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_37), .ScanIn(nScanOut2022), .ScanOut(nScanOut2021), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2022 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_38), .ScanIn(nScanOut2023), .ScanOut(nScanOut2022), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2023 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_39), .ScanIn(nScanOut2024), .ScanOut(nScanOut2023), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2024 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_40), .ScanIn(nScanOut2025), .ScanOut(nScanOut2024), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2025 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_41), .ScanIn(nScanOut2026), .ScanOut(nScanOut2025), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2026 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_42), .ScanIn(nScanOut2027), .ScanOut(nScanOut2026), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2027 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_43), .ScanIn(nScanOut2028), .ScanOut(nScanOut2027), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2028 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_44), .ScanIn(nScanOut2029), .ScanOut(nScanOut2028), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2029 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_45), .ScanIn(nScanOut2030), .ScanOut(nScanOut2029), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2030 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_46), .ScanIn(nScanOut2031), .ScanOut(nScanOut2030), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2031 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_47), .ScanIn(nScanOut2032), .ScanOut(nScanOut2031), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2032 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_48), .ScanIn(nScanOut2033), .ScanOut(nScanOut2032), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2033 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_49), .ScanIn(nScanOut2034), .ScanOut(nScanOut2033), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2034 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_50), .ScanIn(nScanOut2035), .ScanOut(nScanOut2034), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2035 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_51), .ScanIn(nScanOut2036), .ScanOut(nScanOut2035), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2036 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_52), .ScanIn(nScanOut2037), .ScanOut(nScanOut2036), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2037 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_53), .ScanIn(nScanOut2038), .ScanOut(nScanOut2037), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2038 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_54), .ScanIn(nScanOut2039), .ScanOut(nScanOut2038), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2039 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_55), .ScanIn(nScanOut2040), .ScanOut(nScanOut2039), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2040 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_56), .ScanIn(nScanOut2041), .ScanOut(nScanOut2040), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2041 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_57), .ScanIn(nScanOut2042), .ScanOut(nScanOut2041), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2042 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_58), .ScanIn(nScanOut2043), .ScanOut(nScanOut2042), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2043 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_59), .ScanIn(nScanOut2044), .ScanOut(nScanOut2043), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2044 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_60), .ScanIn(nScanOut2045), .ScanOut(nScanOut2044), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2045 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_61), .ScanIn(nScanOut2046), .ScanOut(nScanOut2045), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2046 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_62), .ScanIn(nScanOut2047), .ScanOut(nScanOut2046), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2047 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut31_63), .ScanIn(nScanOut2048), .ScanOut(nScanOut2047), .ScanEnable(nScanEnable) );
Jacobi_Control #( 8, 7, 1, 1 ) U_Jacobi_Control ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Enable(nEnable), .ScanId(1'd0), .ScanEnable(nScanEnable), .ScanIn(nScanOut0), .ScanOut(nScanOut2048) );

/*
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
