`define REG_WIDTH 16
`define REG_SIZE 5
`define ADDRESS_WIDTH 4
`define GPIO_PINS 16
`define FIFO_BIT_SIZE 4

`timescale 1ns / 1ps

module fifo (
	clk,
	reset,
	input_data,
	wen,
	ren,
	output_data,
	empty,
	full);

input clk;
input reset;
input [`REG_WIDTH-1:0]input_data;
input ren;
input wen;
output [`REG_WIDTH-1:0]output_data;
reg [`REG_WIDTH-1:0]output_data;
output empty;
reg empty;
output full;
reg full;

// Defines sizes in terms of bits.
parameter MAX_COUNT = 4'b1111;	// FIFO cap.  This is 16 mem spots.

// The FIFO pointers.
reg [`FIFO_BIT_SIZE-1:0]tail;
reg [`FIFO_BIT_SIZE-1:0]head;
reg [`FIFO_BIT_SIZE-1:0]count;

// The actual memory
reg [`REG_WIDTH:0]fifo_memory[0:MAX_COUNT];

// outputdata is registered and gets the value that tail points to RIGHT NOW.  The
// head points to the last read.  Because of overflow the head and tail
// autowrap.
always @(posedge clk)
begin
	if (reset == 1'b1) begin
		output_data <= 16'h0000;
		head <= 0;
		tail <= 0;
		count <= 0;
		full <= 0;
		empty <= 0;
	end
	else
	begin
		// the output
		output_data <= fifo_memory[tail];

		// the input write
		if (wen == 1'b1 && full == 1'b0)
		begin
			fifo_memory[head] <= input_data;
			// move the head down
	        	head <= head + 1;
		end

		// moving the tail on a read
	      	if (ren == 1'b1 && empty == 1'b0) begin
	       		// READ
			tail <= tail + 1;
		end

		// what to do under different read write scenarios
		case ({ren, wen})
			2'b00:
			begin
				count <= count;
			end
			2'b01:
			begin
				// WRITE
				if (count != MAX_COUNT)
				begin
					count <= count + 1;
				end
	      			empty <= 1'b0;
			end
			2'b10:
			begin
				// READ
				if (count != 2'b00)
				begin
					count <= count - 1;
				end
	      			empty <= 1'b0;
			end
			2'b11:
			begin
				// Concurrent read and write.. no change in count
				count <= count;
	      			empty <= 1'b0;
			end
		endcase

		// full and empty signals
	   	if (count == MAX_COUNT)
		begin
			full <= 1'b1;
		end
		else if (count == 0)
		begin
			empty <= 1'b1;
		end
		else
		begin
			full <= 1'b0;
		end
	end
end

endmodule

`timescale 1ns / 1ps

module gpio_port(
	clk,
	reset,
	gpio_pins,
	INT,
	spi_write_int,
	ready,
	read,
	address,
	value_register_input,
	value_register_output,
	value_wen,
	fifo_write,
	fifo_wen);

input clk;
input reset;

/* the pins coming in */
inout [`GPIO_PINS-1:0]gpio_pins;
/* the gpio_ports in out wires.  This is needed to properly deal with the
* two way nature of the ports */
wire [`GPIO_PINS-1:0]gpio_pins_out;
wire [`GPIO_PINS-1:0]gpio_pins_in;

/* for the chip interrupt on reads or keypresses */
output INT;
wire INT;

/* spi_write_int is a signal which tells if a write happens and we need to
* reinitialize the directions and values of the gpio_pins */
input spi_write_int;
/* tells the control that it can initialize the gpio ports */
input ready;

/* the access pins to the register file */
input [`REG_WIDTH-1:0] read;
output [`ADDRESS_WIDTH-1:0] address;
reg [`ADDRESS_WIDTH-1:0] address;

/* access to the register files value register.  We get direct access since
* it is heavily used */
input [`REG_WIDTH-1:0]value_register_input;
output [`REG_WIDTH-1:0]value_register_output;
wire [`REG_WIDTH-1:0]value_register_output;
output value_wen;
wire value_wen;

/* init direction is the initial state to send out all Zs on the gpios */
reg init_direction;

reg [`GPIO_PINS-1:0]control_register;
/* the register indicating which reading pins interrupt */
reg [`GPIO_PINS-1:0]interrupt_register;
/* the register containing the direction of each gpio_pin.
* 1 = input/reads, 0 = output/writes */
reg [`GPIO_PINS-1:0]direction_register;
/* the values for the right and read registers */
reg [`GPIO_PINS-1:0]value_register;
/* the register for directions of pins in keypad mode */
wire [`GPIO_PINS-1:0]mask_keypad_dir_register;
/* the pins in the keypad that are dedicate for each row and collumn */
wire [`GPIO_PINS-1:0]mask_column_bits; // collumns send out signals
wire [`GPIO_PINS-1:0]mask_row_bits; // rows are read

/* control signals to the two different units of gpio behaviour */
reg gpio_ctrl_ready;
reg keypad_ready;
// this is the interrupt signal generated by the non-keypad pins...
wire gpio_ctrl_interrupt;
wire keypad_interrupt;

/* control of when to write keypresses to the fifo */
output fifo_wen;
wire fifo_wen;
output [`REG_WIDTH-1:0]fifo_write;
wire [`REG_WIDTH-1:0]fifo_write;

/* the output from the keypad controller */
wire [`GPIO_PINS-1:0]keypad_controller_out;

parameter STATE_SIZE=7;
parameter RESET =							7'b0000001, // 01
			INIT =	 					7'b0000010, // 02
			SET_CONTROL_REGISTER =				7'b0000100, // 04
			SET_INT_REGISTER = 				7'b0001000, // 08
			SET_DIRECTION_REGISTER_AND_VALUE_REGISTER = 	7'b0010000, // 10
			NORMAL_OPERATION = 				7'b1000000; // 12

reg [STATE_SIZE-1:0]state;
reg [STATE_SIZE-1:0]next_state;

// module for the keypad controller
keypad_controller kc(
	.clk(clk),
	.reset(reset),
	.gpio_pins_in(gpio_pins_in),
	.keypad_controller_out(keypad_controller_out),
	.row_mask(mask_row_bits),
	.column_mask(mask_column_bits),
	.control_register(control_register),
	.ready(keypad_ready),
	.interrupt(keypad_interrupt),
	.fifo_out(fifo_write),
	.fifo_wen(fifo_wen));

// the controller for the pins in non-keypad mode
gpio_read_pins read_controller(
	.clk(clk),
	.reset(reset),
	.gpio_pins_in(gpio_pins_in),
	.read_mask(direction_register),
	.interrupt_mask(interrupt_register),
	.ready(gpio_ctrl_ready),
	.interrupt(gpio_ctrl_interrupt),
	.value_register_input(value_register_input),
	.value_register_output(value_register_output),
	.value_wen(value_wen));

// figure out the pins that are dedicated for keypad
turn_on_ports pins_used_by_keypad1(control_register[3:0]+{2'b00,control_register[6:4]}, mask_keypad_dir_register);
// figure out the keypad row pins
turn_on_ports pins_used_by_keypad2({1'b0, control_register[3:0]}, mask_row_bits);
// figure out the keypad collumn pins
assign mask_column_bits = mask_keypad_dir_register & ~mask_row_bits;

// simple interrupt behaviour since we just or them
assign INT = gpio_ctrl_interrupt | keypad_interrupt;

// always write out on these pins.  The direction register masks out non writing bis
assign gpio_pins_out = (value_register & ~mask_keypad_dir_register) | (keypad_controller_out & mask_keypad_dir_register);

// mask for the output pins
assign gpio_pins[0] = (init_direction && !direction_register [0]) ? gpio_pins_out[0] : 1'bz;
assign gpio_pins[1] = (init_direction && !direction_register [1]) ? gpio_pins_out[1] : 1'bz;
assign gpio_pins[2] = (init_direction && !direction_register [2]) ? gpio_pins_out[2] : 1'bz;
assign gpio_pins[3] = (init_direction && !direction_register [3]) ? gpio_pins_out[3] : 1'bz;
assign gpio_pins[4] = (init_direction && !direction_register [4]) ? gpio_pins_out[4] : 1'bz;
assign gpio_pins[5] = (init_direction && !direction_register [5]) ? gpio_pins_out[5] : 1'bz;
assign gpio_pins[6] = (init_direction && !direction_register [6]) ? gpio_pins_out[6] : 1'bz;
assign gpio_pins[7] = (init_direction && !direction_register [7]) ? gpio_pins_out[7] : 1'bz;
assign gpio_pins[8] = (init_direction && !direction_register [8]) ? gpio_pins_out[8] : 1'bz;
assign gpio_pins[9] = (init_direction && !direction_register [9]) ? gpio_pins_out[9] : 1'bz;
assign gpio_pins[10] = (init_direction && !direction_register [10]) ? gpio_pins_out[10] : 1'bz;
assign gpio_pins[11] = (init_direction && !direction_register [11]) ? gpio_pins_out[11] : 1'bz;
assign gpio_pins[12] = (init_direction && !direction_register [12]) ? gpio_pins_out[12] : 1'bz;
assign gpio_pins[13] = (init_direction && !direction_register [13]) ? gpio_pins_out[13] : 1'bz;
assign gpio_pins[14] = (init_direction && !direction_register [14]) ? gpio_pins_out[14] : 1'bz;
assign gpio_pins[15] = (init_direction && !direction_register [15]) ? gpio_pins_out[15] : 1'bz;

// mask for the input pins
assign gpio_pins_in[0] = (init_direction && direction_register [0]) ? gpio_pins[0] : 1'bz;
assign gpio_pins_in[1] = (init_direction && direction_register [1]) ? gpio_pins[1] : 1'bz;
assign gpio_pins_in[2] = (init_direction && direction_register [2]) ? gpio_pins[2] : 1'bz;
assign gpio_pins_in[3] = (init_direction && direction_register [3]) ? gpio_pins[3] : 1'bz;
assign gpio_pins_in[4] = (init_direction && direction_register [4]) ? gpio_pins[4] : 1'bz;
assign gpio_pins_in[5] = (init_direction && direction_register [5]) ? gpio_pins[5] : 1'bz;
assign gpio_pins_in[6] = (init_direction && direction_register [6]) ? gpio_pins[6] : 1'bz;
assign gpio_pins_in[7] = (init_direction && direction_register [7]) ? gpio_pins[7] : 1'bz;
assign gpio_pins_in[8] = (init_direction && direction_register [8]) ? gpio_pins[8] : 1'bz;
assign gpio_pins_in[9] = (init_direction && direction_register [9]) ? gpio_pins[9] : 1'bz;
assign gpio_pins_in[10] = (init_direction && direction_register [10]) ? gpio_pins[10] : 1'bz;
assign gpio_pins_in[11] = (init_direction && direction_register [11]) ? gpio_pins[11] : 1'bz;
assign gpio_pins_in[12] = (init_direction && direction_register [12]) ? gpio_pins[12] : 1'bz;
assign gpio_pins_in[13] = (init_direction && direction_register [13]) ? gpio_pins[13] : 1'bz;
assign gpio_pins_in[14] = (init_direction && direction_register [14]) ? gpio_pins[14] : 1'bz;
assign gpio_pins_in[15] = (init_direction && direction_register [15]) ? gpio_pins[15] : 1'bz;

always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		init_direction <= 1'b0; // makesure nothing is written out or accepted until the first initlization sequence is done
		direction_register <= 0;
		interrupt_register <= 0;
		value_register <= 0;
		control_register <= 0;
		gpio_ctrl_ready <= 1'b0; // this controls the reading interrupt and writing control
		address <= 0;
		keypad_ready <= 1'b0; // this controls the keypad reader
	end
	else
	begin
		case (state)
			INIT:
			begin
				/* read control register */
				address <= 0;
			end
			SET_CONTROL_REGISTER:
			begin
				/* read interrupt register */
				address <= 1;
				control_register <= read;
			end
			SET_INT_REGISTER:
			begin
				/* read direction register */
				address <= 2;
				interrupt_register <= read;
			end
			SET_DIRECTION_REGISTER_AND_VALUE_REGISTER:
			begin
				direction_register <= ((read & ~mask_keypad_dir_register) | mask_row_bits); // first part picks reads not in use by keypda.  Last or picks the row bits which will be reads
				/* read value register - can read right away since we get port directly */
				value_register <= (value_register_input & ~direction_register); // only put in write bits
			end
			NORMAL_OPERATION:
			begin
				init_direction <= 1'b1;
				gpio_ctrl_ready <= 1'b1;
				keypad_ready <= 1'b1;
			end
			default:
			begin
			end
		endcase

	end
end

/* Combinational state machine */
always @(state or ready or spi_write_int)
begin
	next_state = 0;
	case (state)
		RESET:
		begin
			if (ready == 1'b1)
			begin
				next_state = INIT;
			end
			else
			begin
				next_state = RESET;
			end
		end
		INIT:
		begin
			next_state = SET_CONTROL_REGISTER;
		end
		SET_CONTROL_REGISTER:
		begin
			if (spi_write_int == 1'b1)
			begin
				next_state = INIT;
			end
			else
			begin
				next_state = SET_INT_REGISTER;
			end
		end
		SET_INT_REGISTER:
		begin
			if (spi_write_int == 1'b1)
			begin
				next_state = INIT;
			end
			else
			begin
				next_state = SET_DIRECTION_REGISTER_AND_VALUE_REGISTER;
			end
		end
		SET_DIRECTION_REGISTER_AND_VALUE_REGISTER:
		begin
			if (spi_write_int == 1'b1)
			begin
				next_state = INIT;
			end
			else
			begin
				next_state = NORMAL_OPERATION;
			end
		end
		NORMAL_OPERATION:
		begin
			if (spi_write_int == 1'b1)
			begin
				next_state = INIT;
			end
			else
			begin
				next_state = NORMAL_OPERATION;
			end
		end
		default:
		begin
			next_state = INIT;
		end
	endcase
end

/* sequential state changes */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		state <= RESET;
		next_state <= RESET;
	end
	else
	begin
		state <= next_state;
	end
end

endmodule

`timescale 1ns / 1ps

module gpio_read_pins(
	clk,
	reset,
	gpio_pins_in,
	read_mask,
	interrupt_mask,
	ready,
	interrupt,
	value_register_input,
	value_register_output,
	value_wen);

input clk;
input reset;

/* the gpio_pins input is the only things needed to be handled...when they
* change */
input [`GPIO_PINS-1:0]gpio_pins_in;
/* masks for what is to be read and interrupted on */
input [`GPIO_PINS-1:0]read_mask;
input [`GPIO_PINS-1:0]interrupt_mask;
/* signal to indicate when this device can begin normal operation */
input ready;

// the pin we send interrupts on for 1 cycle ... the gpio then decides which interrupt to send
output interrupt;
reg interrupt;

// direct access to writing of value register in reg file
input [`REG_WIDTH-1:0]value_register_input;
output [`REG_WIDTH-1:0]value_register_output;
wire [`REG_WIDTH-1:0]value_register_output;
output value_wen;
reg value_wen;

/* registers and wires to handle logic for changes on these pins */
reg [`GPIO_PINS-1:0]last_in_value;
reg [`GPIO_PINS-1:0]last_in_value_int;
wire [`GPIO_PINS-1:0]in_value;
wire [`GPIO_PINS-1:0]in_value_int;
wire [`GPIO_PINS-1:0]change;
wire [`GPIO_PINS-1:0]change_int;

parameter STATE_SIZE=4;
parameter RESET =			4'b0001,
			IDLE =	 	4'b0010,
			INTERRUPT = 	4'b0100,
			UPDATE = 	4'b1000;

reg [STATE_SIZE-1:0]state;
reg [STATE_SIZE-1:0]next_state;

// always have the write going out...needs to be activated with the value_wen
assign value_register_output = (value_register_input & ~read_mask) | (gpio_pins_in & read_mask);
// mask in the reads that and the reads that should be interrupted
assign in_value = gpio_pins_in & read_mask;
assign in_value_int = gpio_pins_in & read_mask & interrupt_mask;
// bitwise xor to see if there is a change
assign change = in_value ^ last_in_value;
assign change_int = in_value_int ^ last_in_value_int;

always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		interrupt <= 1'b0;
		value_wen <= 1'b0;
	end
	else
	begin
		case (state)
			IDLE:
			begin
				interrupt <= 1'b0;
				value_wen <= 1'b0;
			end
			INTERRUPT:
			begin
				interrupt <= 1'b1; // interrupt since changed on interrupt pin
				value_wen <= 1'b1; // write value since changed
			end
			UPDATE:
			begin
				interrupt <= 1'b0;
				value_wen <= 1'b1; // write value since changed
			end
		endcase

	end
end

/* Combinational state machine */
always @(state or ready or change or change_int)
begin
	next_state = 0;
	case (state)
		RESET:
		begin
			if (ready == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = RESET;
			end
		end
		IDLE:
		begin
			if (change_int != 0)
			begin
				next_state = INTERRUPT;
			end
			else if (change != 0)
			begin
				next_state = UPDATE;
			end
			else
			begin
				next_state = IDLE;
			end
		end
		INTERRUPT:
		begin
			next_state = IDLE;
		end
		UPDATE:
		begin
			next_state = IDLE;
		end
		default:
		begin
			next_state = RESET;
		end
	endcase
end

/* sequential state changes */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		state <= RESET;
		next_state <= RESET;
		last_in_value_int <= 0;
		last_in_value <= 0;
	end
	else
	begin
		state <= next_state;
		// keep a record so we can figure out changes
		last_in_value_int <= in_value_int;
		last_in_value <= in_value;
	end
end

endmodule

`timescale 1ns / 1ps

module io_expander(
	clk,
	reset,
	SCLK,
	SI,
	SO,
	SS,
	INT,
	gpio_pins);

input clk;
input reset;

/* SPI pins */
input SCLK;
input SI;
input SS;
output SO;
wire SO;

/* the general purpose io pins */
inout [`GPIO_PINS-1:0]gpio_pins;

/* interrupt signal */
output INT;
wire INT;

/* access wires to the register file */
wire [`REG_WIDTH-1:0] read;
wire [`REG_WIDTH-1:0] write;
wire [`ADDRESS_WIDTH-1:0] address_regfile;
wire [`ADDRESS_WIDTH-1:0] address_gpio;
wire [`ADDRESS_WIDTH-1:0] address_spi;
wire wen;

/* bit to tell the device when it has all the registers properly programmed
* and can operate */
wire ready_bit;

/* bit to tell if there is a new programming of the chip and we need to
* reset the keypad and gpio control structures */
reg spi_write_int;
/* a bit that tells the gpio when it can operate */
reg gpio_ready;

/* wires for direct access of the value register in the register file */
wire [`REG_WIDTH-1:0] value_register_in;
wire [`REG_WIDTH-1:0] value_register_out;
wire value_wen;

/* fifo access pins.  Keypad writes, SPI reads on address 5 */
wire fifo_ren;
wire [`REG_WIDTH-1:0]fifo_out;
wire fifo_empty;
wire fifo_wen;
wire [`REG_WIDTH-1:0]fifo_in;
wire fifo_full;

parameter STATE_SIZE=4;
parameter RESET =			4'b0001,
			IDLE =	 	4'b0010;
reg [STATE_SIZE-1:0]state;
reg [STATE_SIZE-1:0]next_state;

/* Register file:
* 0 Control Register
* 1 Interrupt Register A * 2 Interrupt Register B
* 2 Direction Register A * 4 Direction Register B
* 3 Value Register A * 6 Value Register B
* 4 Interrupt Type Register // Not used in this design
* 5 FIFO head */
register_file regfile(
	.clk(clk),
	.reset(reset),
	.out(read),
	.in(write),
	.address(address_regfile),
	.wen(wen),
	.value_register_in(value_register_out),
	.value_register_out(value_register_in),
	.value_wen(value_wen),
	.ready_bit(ready_bit));

spi_interface spi(
	.clk(clk),
	.reset(reset),
	.SCLK(SCLK),
	.SI(SI),
	.SO(SO),
	.SS(SS),
	.read(read),
	.write(write),
	.address(address_spi),
	.wen(wen),
	.fifo_top_entry(fifo_out),
	.fifo_ren(fifo_ren),
	.fifo_empty(fifo_empty));

gpio_port gp(
	.clk(clk),
	.reset(reset),
	.gpio_pins(gpio_pins),
	.INT(INT),
	.spi_write_int(spi_write_int),
	.ready(gpio_ready),
	.read(read),
	.address(address_gpio),
	.value_register_input(value_register_in),
	.value_register_output(value_register_out),
	.value_wen(value_wen),
	.fifo_write(fifo_in),
	.fifo_wen(fifo_wen));

fifo fifo_for_keypresses (
	.clk(clk),
	.reset(reset),
	.input_data(fifo_in),
	.wen(fifo_wen),
	.ren(fifo_ren),
	.output_data(fifo_out),
	.empty(fifo_empty),
	.full(fifo_full));

/* another poor way of accessing memory.  If both try to access at the same
* time we'll have trouble */
assign address_regfile = address_spi | address_gpio;

always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		gpio_ready <= 1'b0;
	end
	else
	begin
		case (state)
			IDLE:
			begin
				gpio_ready <= 1'b1;
			end
		endcase

	end
end

/* Combinational state machine */
always @(state or ready_bit)
begin
	next_state = 0;
	case (state)
		RESET:
		begin
			if (ready_bit == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = RESET;
			end
		end
		IDLE:
		begin
			next_state = IDLE;
		end
		default:
		begin
			next_state = RESET;
		end
	endcase
end

/* sequential state changes */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		state <= RESET;
		next_state <= RESET;
	end
	else
	begin
		state <= next_state;
	end
end

endmodule

`timescale 1ns / 1ps

module keygrid_4x4 (
	presses,
	column_ins,
	row_outs);

// This helps testing of a 4x4 keypad by sending signals out based on the
// incoming high signals.  The theoretical keypad is as below
/*     0  1  2  3
*   -------------
*   0| 0  1  2  3
*   1| 4  5  6  7
*   2| 8  9  10 11
*   3| 12 13 14 15
*/
input [15:0]presses;
input [3:0]column_ins;
output [3:0]row_outs;
wire [3:0]row_outs;

assign row_outs[0] = ((presses[0] == 1'b1 && column_ins[0] == 1'b1) || (presses[1] == 1'b1 && column_ins[1] == 1'b1) || (presses[2] == 1'b1 && column_ins[2] == 1'b1) || (presses[3] == 1'b1 && column_ins[3] == 1'b1)) ? 1'b1 : 1'b0;
assign row_outs[1] = ((presses[4] == 1'b1 && column_ins[0] == 1'b1) || (presses[5] == 1'b1 && column_ins[1] == 1'b1) || (presses[6] == 1'b1 && column_ins[2] == 1'b1) || (presses[7] == 1'b1 && column_ins[3] == 1'b1)) ? 1'b1 : 1'b0;
assign row_outs[2] = ((presses[8] == 1'b1 && column_ins[0] == 1'b1) || (presses[9] == 1'b1 && column_ins[1] == 1'b1) || (presses[10] == 1'b1 && column_ins[2] == 1'b1) || (presses[11] == 1'b1 && column_ins[3] == 1'b1)) ? 1'b1 : 1'b0;
assign row_outs[3] = ((presses[12] == 1'b1 && column_ins[0] == 1'b1) || (presses[13] == 1'b1 && column_ins[1] == 1'b1) || (presses[14] == 1'b1 && column_ins[2] == 1'b1) || (presses[15] == 1'b1 && column_ins[3] == 1'b1)) ? 1'b1 : 1'b0;

endmodule


`timescale 1ns / 1ps

module keypad_controller(
	clk,
	reset,
	gpio_pins_in,
	keypad_controller_out,
	row_mask,
	column_mask,
	control_register,
	ready,
	interrupt,
	fifo_out,
	fifo_wen);

input clk;
input reset;

/* gpio pins in */
input [`GPIO_PINS-1:0]gpio_pins_in;
/* what the keypad controller will send out in terms of signals */
output [`GPIO_PINS-1:0]keypad_controller_out;
wire [`GPIO_PINS-1:0]keypad_controller_out;

// the masks for which pins do what
input [`GPIO_PINS-1:0]row_mask;
input [`GPIO_PINS-1:0]column_mask;

// control register for which pins are what in the keypad
input [`GPIO_PINS-1:0]control_register;

// the signal that tells the keypad controller to start
input ready;

// the pin we send interrupts on for 1 cycle ... the gpio then decides which interrupt to send
output interrupt;
reg interrupt;

// direct access to writing of value register in reg file
output [`REG_WIDTH-1:0]fifo_out;
reg [`REG_WIDTH-1:0]fifo_out;
output fifo_wen;
reg fifo_wen;

// pins that are supposed to be active as polling pins
wire [`GPIO_PINS-1:0]active_poll_pins;
// counters as we go through the polling
reg [3:0]row_counter;
reg [3:0]column_counter;

// records the changes and compares against the current signal.  last
// keypress is for storing a keypress before polling
reg [`GPIO_PINS-1:0]last_in_value;
reg [`GPIO_PINS-1:0]last_keypress;
wire [`GPIO_PINS-1:0]change;
wire [`REG_WIDTH-1:0]in_value;

parameter STATE_SIZE=6;
parameter RESET =				6'b000001,
			IDLE =			6'b000010,
			CHANGE = 		6'b000100,
			POLL_NEXT_COLUMN =	6'b001000,
			POLL_NEXT_ROWS = 	6'b010000,
			DONE_POLL = 		6'b100000;

reg [STATE_SIZE-1:0]state;
reg [STATE_SIZE-1:0]next_state;

// depending on counter returns an active vector for polling
turn_on_poll_pins topp({1'b0, column_counter}, active_poll_pins);

// mask in the reads that and the reads that should be interrupted
assign /*in_value*/in_value = gpio_pins_in & row_mask;
// bitwise xor to see if there is a change
assign change = in_value ^ last_in_value;
//      		          the non-keypad value   the collumn output pins masked
assign keypad_controller_out = (active_poll_pins & (column_mask & ~row_mask));

always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		interrupt <= 1'b0;
		fifo_wen <= 1'b0;
		column_counter <= 0; // set to value the number of columns
		last_keypress <= 0;
		fifo_out <= 0;
	end
	else
	begin
		case (state)
			IDLE:
			begin
				interrupt <= 1'b0;
				column_counter <= 0; // set to value the number of columns
			end
			CHANGE:
			begin
				last_keypress <= in_value; // record the keypress so we can restore last_in_value after polling keypad
				column_counter <= control_register[3:0]; // start at the number of rows since those low pins (rows) are for reading
				row_counter <= 0; // set to value of the number of rows
			end
			POLL_NEXT_COLUMN:
			begin
				// increase the counter to set a different pin
				column_counter <= column_counter + 1; // this increase will also change the polling output pin
				row_counter <= 0;
				fifo_wen <= 1'b0;
			end
			POLL_NEXT_ROWS:
			begin
				row_counter <= row_counter + 1;
				if (in_value[row_counter] != 0)
				begin
					/* if there is a value then we've found a keypress so write to the fifo */
					fifo_wen <= 1'b1;
					fifo_out <= {column_counter-control_register[6:4],row_counter};
				end
				else
				begin
					fifo_wen <= 1'b0;
					fifo_out <= 0;
				end
			end
			DONE_POLL:
			begin
				/* after a poll send an interrupt */
				interrupt <= 1'b1;
				/* turn off the fifo wren just in case it was on */
				fifo_wen <= 1'b0;
			end
		endcase
	end
end

/* Combinational state machine */
always @(state or ready or change or column_counter or row_counter)
begin
	next_state = 0;
	case (state)
		RESET:
		begin
			if (ready == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = RESET;
			end
		end
		IDLE:
		begin
			if (ready == 1'b0)
			begin
				next_state = RESET;
			end
			else if (change != 0)
			begin
				next_state = CHANGE;
			end
			else
			begin
				next_state = IDLE;
			end
		end
		CHANGE:
		begin
			if (ready == 1'b0)
			begin
				next_state = RESET;
			end
			else
			begin
				next_state = POLL_NEXT_COLUMN;
			end
		end
		POLL_NEXT_COLUMN:
		begin
			if (ready == 1'b0)
			begin
				next_state = RESET;
			end
			else if (column_counter == control_register[6:4]+control_register[6:4])
			begin
				next_state = DONE_POLL;
			end
			else
			begin
				next_state = POLL_NEXT_ROWS;
			end
		end
		POLL_NEXT_ROWS:
		begin
			if (ready == 1'b0)
			begin
				next_state = RESET;
			end
			else if (row_counter == control_register[3:0]-1)
			begin
				next_state = POLL_NEXT_COLUMN;
			end
			else
			begin
				next_state = POLL_NEXT_ROWS;
			end
		end
		DONE_POLL:
		begin
			if (ready == 1'b0)
			begin
				next_state = RESET;
			end
			else
			begin
				next_state = IDLE;
			end
		end
		default:
		begin
			next_state = RESET;
		end
	endcase
end

/* sequential state changes */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		state <= RESET;
		next_state <= RESET;
		last_in_value <= in_value;
	end
	else
	begin
		state <= next_state;
		// keep a record so we can figure out changes
		if (state == IDLE)
		begin
			// update the last in_value with the last keypress
			last_in_value <= last_keypress;
		end
		else
		begin
			/* otherwise record old state to check for changes */
			last_in_value <= in_value;
		end
	end
end

endmodule

`timescale 1ns / 1ps

module register_file(clk, reset, out, in, address, wen, value_register_in, value_register_out, value_wen, ready_bit);

/* Register file:
* 0 Control Register
* 1 Interrupt Register A * 2 Interrupt Register B
* 2 Direction Register A * 4 Direction Register B
* 3 Value Register A * 6 Value Register B
* 4 Interrupt Type Register
* 5 is fifo head, but not part of register file */

input clk;
input reset;
output [`REG_WIDTH-1:0] out;
wire [`REG_WIDTH-1:0] out;
input [`REG_WIDTH-1:0] in;
input [`ADDRESS_WIDTH-1:0] address;
input wen;

/* specialised direct connections so other parts of the circuit can
* directly access the value register */
input [`REG_WIDTH-1:0] value_register_in;
input value_wen;
output [`REG_WIDTH-1:0] value_register_out;
wire [`REG_WIDTH-1:0] value_register_out;

/* special bit that is set in register when all the data is in from the
* control register to setup the device operation */
output ready_bit;
wire ready_bit;

/* register file */
reg [`REG_WIDTH-1:0] registers [`REG_SIZE-1:0];

/* always send out address 3 */
assign value_register_out = registers[3];
/* link to the ready bit in the control register */
assign ready_bit = registers[0][8];
/* the output of the register file */
assign out = registers[address];

always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
	end
	else
	begin
		if (wen == 1'b1)
		begin
			registers[address] <= in;
		end

		if (value_wen == 1'b1)
		begin
			registers[3] <= value_register_in;
		end
	end
end

endmodule



`timescale 1ns / 1ps

module spi_interface(
	clk,
	reset,
	SCLK,
	SI,
	SO,
	SS,
	read,
	write,
	address,
	wen,
	fifo_top_entry,
	fifo_ren,
	fifo_empty);

input clk;
input reset;

/* access to the register file */
input [`REG_WIDTH-1:0] read;
output [`REG_WIDTH-1:0] write;
output [`ADDRESS_WIDTH-1:0] address;
reg [`ADDRESS_WIDTH-1:0] address;
output wen;
reg wen;
wire [`REG_WIDTH-1:0] write;

/* the SPI pins */
input SCLK;
input SI;
output SO;
reg SO;
input SS;

/* counters to count SCLK and packets */
reg [4:0]clock_counter;
reg [1:0]packets;

/* the actual read register */
reg [15:0]spi_read_register;

/* the fifo read port */
input [`REG_WIDTH-1:0] fifo_top_entry;
output fifo_ren;
reg fifo_ren;
input fifo_empty;

parameter STATE_SIZE=11;
parameter IDLE = 									11'b00000000001,//001
			INPUT_READ = 							11'b00000000010,//002
			INPUT_READ_CLOCK_HIGH_COUNT = 	11'b00000000100,//004
			INPUT_READ_CLOCK_HIGH = 			11'b00000001000,//008
			INPUT_READ_CLOCK_LOW_SAMPLE = 	11'b00000010000,//010
			INPUT_READ_CLOCK_LOW = 				11'b00000100000,//020
			OUTPUT_READ_CLOCK_HIGH_COUNT = 	11'b00100000000,//100
			OUTPUT_READ_CLOCK_HIGH = 			11'b01000000000,//200
			OUTPUT_READ_CLOCK_LOW =			 	11'b10000000000;//400

reg [STATE_SIZE-1:0]state;
reg [STATE_SIZE-1:0]next_state;

/* the write always goes out */
assign write = spi_read_register;

/* output logic */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		clock_counter <= 0;
		SO <= 1'bx;
		spi_read_register <= 0;
		packets <= 0;
		fifo_ren <= 1'b0;
	end
	else
	begin
		case (state)
			IDLE:
			begin
				wen <= 1'b0;
				SO <= 1'bx;
				spi_read_register <= 0;
				packets <= 0;
				fifo_ren <= 1'b0;
			end
			INPUT_READ:
			begin
				// in read mode reset the clock counter
				clock_counter <= 0;
			end
			INPUT_READ_CLOCK_HIGH_COUNT:
			begin
				// found high bit so count next clock
				clock_counter <= clock_counter + 1;
			end
			INPUT_READ_CLOCK_HIGH:
			begin
			end
			INPUT_READ_CLOCK_LOW_SAMPLE:
			begin
				// record the value in the spi_read_register
				spi_read_register[clock_counter-1] <= SI;
			end
			INPUT_READ_CLOCK_LOW:
			begin
				if ((((clock_counter == 8) && (packets == 0)) || ((clock_counter == 16) && (packets == 1))) && (SS == 1'b0))
				begin
					if ((spi_read_register[0] == 1'b1) && (packets == 0)) // read 16 bits
					begin
						address <= spi_read_register[4:1];
						spi_read_register <= 0;
						wen <= 1'b0;
						clock_counter <= 0;
						packets <= packets + 1;
					end
					else // 0 = write
					begin
						clock_counter <= 0;
						if (packets == 0)
						begin
							// set up the writing
							address <= spi_read_register[4:1];
							spi_read_register <= 0;
							packets <= packets + 1;
						end
						else
						begin
							// write the second read value
							wen <= 1'b1;
						end
					end
				end
			end
			OUTPUT_READ_CLOCK_HIGH_COUNT:
			begin
				// read is actaully an output since the
				// external world wants to read a register
				//
				// count the clocks
				clock_counter <= clock_counter + 1;
			end
			OUTPUT_READ_CLOCK_HIGH:
			begin
				if (address == 5) // if we're reading from the fifo of keypresses
				begin
					if (fifo_empty == 1'b0)
					begin
						SO <= fifo_top_entry[clock_counter-1];
					end
					else
					begin
						SO <= 0;
					end
				end
				else
				begin
					// sendout the read register form the file
					SO <= read[clock_counter-1];
				end
			end
			OUTPUT_READ_CLOCK_LOW:
			begin
				if ((clock_counter == 16) && (SS == 1'b0))
				begin
					// if we count the last bit
					if (address == 5) // if we're reading from the fifo of keypresses
					begin
						if (fifo_empty == 1'b0)
						begin
							fifo_ren <= 1'b1; // move the fifo to the next item
						end
					end
				end
			end
			default:
			begin
			end
		endcase
	end
end

/* Combinational state machine */
always @(state or SCLK or SS or clock_counter or spi_read_register or packets)
begin
	next_state = 0;
	case (state)
		IDLE:
		begin
			if ((SCLK == 1'b1) && (SS == 1'b0)) // SS is active low
			begin
				next_state = INPUT_READ;
			end
			else
			begin
				next_state = IDLE;
			end
		end
		INPUT_READ:
		begin
			if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = INPUT_READ_CLOCK_HIGH_COUNT;
			end
		end
		INPUT_READ_CLOCK_HIGH_COUNT:
		begin
			// Waiting for clock to go low so we can read bit and count bits read
			if ((SCLK == 1'b0) && (SS == 1'b0))
			begin
				next_state = INPUT_READ_CLOCK_LOW_SAMPLE;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = INPUT_READ_CLOCK_HIGH;
			end
		end
		INPUT_READ_CLOCK_HIGH:
		begin
			// Waiting for clock to go low so we can read bit and count bits read
			if ((SCLK == 1'b0) && (SS == 1'b0))
			begin
				next_state = INPUT_READ_CLOCK_LOW_SAMPLE;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = INPUT_READ_CLOCK_HIGH;
			end
		end
		INPUT_READ_CLOCK_LOW_SAMPLE:
		begin
			// Waiting for clock to go high
			if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = INPUT_READ_CLOCK_LOW;
			end
		end
		INPUT_READ_CLOCK_LOW:
		begin
			// Waiting for clock to go high
			if ((((clock_counter == 8) && (packets == 0)) ||  ((clock_counter == 16) && (packets == 1))) && (SS == 1'b0))
			begin
				if ((spi_read_register[0] == 1'b1) && (packets == 0)) // read
				begin
					next_state = OUTPUT_READ_CLOCK_LOW;
				end
				else if (packets == 0) // 0 = write
				begin
					next_state = INPUT_READ;
				end
				else
				begin
					next_state = IDLE;
				end
			end
			else if ((SCLK == 1'b1) && (SS == 1'b0))
			begin
				next_state = INPUT_READ_CLOCK_HIGH_COUNT;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = INPUT_READ_CLOCK_LOW;
			end
		end
		OUTPUT_READ_CLOCK_HIGH_COUNT:
		begin
			// Waiting for clock to go low so we can read bit and count bits read
			if ((SCLK == 1'b0) && (SS == 1'b0))
			begin
				next_state = OUTPUT_READ_CLOCK_LOW;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = OUTPUT_READ_CLOCK_HIGH;
			end
		end
		OUTPUT_READ_CLOCK_HIGH:
		begin
			// Waiting for clock to go low so we can read bit and count bits read
			if ((SCLK == 1'b0) && (SS == 1'b0))
			begin
				next_state = OUTPUT_READ_CLOCK_LOW;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = OUTPUT_READ_CLOCK_HIGH;
			end
		end
		OUTPUT_READ_CLOCK_LOW:
		begin
			// Waiting for clock to go high
			if ((clock_counter == 16) && (SS == 1'b0))
			begin
				next_state = IDLE;
			end
			else if ((SCLK == 1'b1) && (SS == 1'b0))
			begin
				next_state = OUTPUT_READ_CLOCK_HIGH_COUNT;
			end
			else if (SS == 1'b1)
			begin
				next_state = IDLE;
			end
			else
			begin
				next_state = OUTPUT_READ_CLOCK_LOW;
			end
		end
		default:
		begin
			next_state = IDLE;
		end
	endcase
end

/* sequential state changes */
always @(posedge clk or posedge reset)
begin
	if (reset == 1'b1)
	begin
		state <= IDLE;
		next_state <= IDLE;
	end
	else
	begin
		state <= next_state;
	end
end

endmodule

`timescale 1ns / 1ps

module turn_on_ports(integers, ones_on);

// simple module that turns on each pin based on the integer value coming in
input [4:0]integers;

output [15:0]ones_on;
wire [15:0]ones_on;

assign ones_on[0] = (integers >= 1) ? 1'b1 : 1'b0;
assign ones_on[1] = (integers >= 2) ? 1'b1 : 1'b0;
assign ones_on[2] = (integers >= 3) ? 1'b1 : 1'b0;
assign ones_on[3] = (integers >= 4) ? 1'b1 : 1'b0;
assign ones_on[4] = (integers >= 5) ? 1'b1 : 1'b0;
assign ones_on[5] = (integers >= 6) ? 1'b1 : 1'b0;
assign ones_on[6] = (integers >= 7) ? 1'b1 : 1'b0;
assign ones_on[7] = (integers >= 8) ? 1'b1 : 1'b0;
assign ones_on[8] = (integers >= 9) ? 1'b1 : 1'b0;
assign ones_on[9] = (integers >= 10) ? 1'b1 : 1'b0;
assign ones_on[10] = (integers >= 11) ? 1'b1 : 1'b0;
assign ones_on[11] = (integers >= 12) ? 1'b1 : 1'b0;
assign ones_on[12] = (integers >= 13) ? 1'b1 : 1'b0;
assign ones_on[13] = (integers >= 14) ? 1'b1 : 1'b0;
assign ones_on[14] = (integers >= 15) ? 1'b1 : 1'b0;
assign ones_on[15] = (integers >= 16) ? 1'b1 : 1'b0;

endmodule

`timescale 1ns / 1ps

module turn_on_poll_pins(integers, ones_on);

// simple module that turns on all pins for 0 otherwise the pin that the
// integer references in the vector
input [4:0]integers;

output [15:0]ones_on;
wire [15:0]ones_on;

assign ones_on[0] = ((integers == 1) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[1] = ((integers == 2) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[2] = ((integers == 3) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[3] = ((integers == 4) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[4] = ((integers == 5) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[5] = ((integers == 6) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[6] = ((integers == 7) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[7] = ((integers == 8) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[8] = ((integers == 9) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[9] = ((integers == 10) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[10] = ((integers == 11) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[11] = ((integers == 12) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[12] = ((integers == 13) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[13] = ((integers == 14) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[14] = ((integers == 15) || (integers == 0)) ? 1'b1 : 1'b0;
assign ones_on[15] = ((integers == 16) || (integers == 0)) ? 1'b1 : 1'b0;

endmodule
