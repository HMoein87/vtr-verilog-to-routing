

/*
 *
 * RAW Benchmark Suite main defines
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/bubblesort/src/library.v,v 1.4 1997/08/09 05:56:59 jbabb Exp $
 *
 * Library for Bubble Sort Benchmark
 *
 * Authors: Elliot Waingold         (elliotw@lcs.mit.edu)
 *          Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 BubbleSort_Node is the basic pairwise element comparator.  It
 outputs the greater of its two inputs to HiOut and the lower of
 the two to LoOut.
 */

module BubbleSort_Node (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
			AIn, BIn, HiOut, LoOut);

   parameter WIDTH = 8;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* local connections */

   input [WIDTH-1:0]		AIn, BIn;
   output [WIDTH-1:0]		HiOut, LoOut;
   wire				Predicate;

   assign Predicate = (AIn > BIn) ? 1 : 0;
   assign HiOut = (Predicate) ? AIn : BIn;
   assign LoOut = (Predicate) ? BIn : AIn;

endmodule


/*
 BubbleSort_Reg is a pipeline/input register that can be written
 to from the host interface as well as from its input wires.  It
 also has an enable input that must be high for it to clock data
 in from the inputs.
 */

module BubbleSort_Reg (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		       ScanIn, ScanOut, ScanEnable,
		       Id, Enable, In, Out);

   parameter			 WIDTH = 8,
				 IDWIDTH = 8,
				 SCAN = 1;

   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;


   /* local connections */

   input [IDWIDTH-1:0]		Id;
   input			Enable;
   input [WIDTH-1:0]		In;
   output [WIDTH-1:0]		Out;
   reg [WIDTH-1:0]		Out;


   /* support reading of the node data value (non-scan only) */

   assign DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out : `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;


   always @(posedge Clk)
      begin


	 /* reset will initialize the register to zero */

	 if (Reset)
	    Out = 0;


	 /* support scan in */

	 else if  (SCAN && ScanEnable)
	    Out = ScanIn[WIDTH-1:0];


	 /* support writing of the node data value (non-scan only) */

	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0] == Id))
	    Out = DataIn[WIDTH-1:0];

	 /* otherwise if enable is high, read in input data */

	 else if (Enable)
	    Out = In;

      end
endmodule


/*
 BubbleSort_Control is the control node.  When a value is written to
 it by the host, it holds the enable high for that number of clock
 periods.
 */

module BubbleSort_Control(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
			  ScanIn, ScanOut, ScanEnable, ScanId,
			  Id, Enable);

   parameter			 CWIDTH=8,
				 IDWIDTH=8,
				 WIDTH=8,
				 SCAN=1;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;
   input [IDWIDTH-1:0]		 ScanId;


   /* local connections */

   input [IDWIDTH-1:0]		 Id;
   output			 Enable;
   reg [CWIDTH-1:0]		 count;
   reg [WIDTH-1:0]		 ScanReg;


   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? count :
         (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;

   /* enable when count is active */

   assign Enable = !(count==0);


   always @(posedge Clk)
      begin


	 /* store current scan output */

	 ScanReg=ScanIn;


	 /* Logic to reset, write, and decrement the counter */

	 if (Reset)
	    count=0;
	 else if (WR && (Addr[IDWIDTH-1:0]==Id))
	    count=DataIn[CWIDTH-1:0];
	 else
	    if(count)
	       count=count-1;
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [31:0] wRegInA0;
wire [31:0] wRegInB0;
wire [31:0] wAIn0;
wire [31:0] wBIn0;
wire [31:0] wRegInA1;
wire [31:0] wRegInB1;
wire [31:0] wAIn1;
wire [31:0] wBIn1;
wire [31:0] wRegInA2;
wire [31:0] wRegInB2;
wire [31:0] wAIn2;
wire [31:0] wBIn2;
wire [31:0] wRegInA3;
wire [31:0] wRegInB3;
wire [31:0] wAIn3;
wire [31:0] wBIn3;
wire [31:0] wRegInA4;
wire [31:0] wRegInB4;
wire [31:0] wAIn4;
wire [31:0] wBIn4;
wire [31:0] wRegInA5;
wire [31:0] wRegInB5;
wire [31:0] wAIn5;
wire [31:0] wBIn5;
wire [31:0] wRegInA6;
wire [31:0] wRegInB6;
wire [31:0] wAIn6;
wire [31:0] wBIn6;
wire [31:0] wRegInA7;
wire [31:0] wRegInB7;
wire [31:0] wAIn7;
wire [31:0] wBIn7;
wire [31:0] wRegInA8;
wire [31:0] wRegInB8;
wire [31:0] wAIn8;
wire [31:0] wBIn8;
wire [31:0] wRegInA9;
wire [31:0] wRegInB9;
wire [31:0] wAIn9;
wire [31:0] wBIn9;
wire [31:0] wRegInA10;
wire [31:0] wRegInB10;
wire [31:0] wAIn10;
wire [31:0] wBIn10;
wire [31:0] wRegInA11;
wire [31:0] wRegInB11;
wire [31:0] wAIn11;
wire [31:0] wBIn11;
wire [31:0] wRegInA12;
wire [31:0] wRegInB12;
wire [31:0] wAIn12;
wire [31:0] wBIn12;
wire [31:0] wRegInA13;
wire [31:0] wRegInB13;
wire [31:0] wAIn13;
wire [31:0] wBIn13;
wire [31:0] wRegInA14;
wire [31:0] wRegInB14;
wire [31:0] wAIn14;
wire [31:0] wBIn14;
wire [31:0] wRegInA15;
wire [31:0] wRegInB15;
wire [31:0] wAIn15;
wire [31:0] wBIn15;
wire [31:0] wRegInA16;
wire [31:0] wRegInB16;
wire [31:0] wAIn16;
wire [31:0] wBIn16;
wire [31:0] wRegInA17;
wire [31:0] wRegInB17;
wire [31:0] wAIn17;
wire [31:0] wBIn17;
wire [31:0] wRegInA18;
wire [31:0] wRegInB18;
wire [31:0] wAIn18;
wire [31:0] wBIn18;
wire [31:0] wRegInA19;
wire [31:0] wRegInB19;
wire [31:0] wAIn19;
wire [31:0] wBIn19;
wire [31:0] wRegInA20;
wire [31:0] wRegInB20;
wire [31:0] wAIn20;
wire [31:0] wBIn20;
wire [31:0] wRegInA21;
wire [31:0] wRegInB21;
wire [31:0] wAIn21;
wire [31:0] wBIn21;
wire [31:0] wRegInA22;
wire [31:0] wRegInB22;
wire [31:0] wAIn22;
wire [31:0] wBIn22;
wire [31:0] wRegInA23;
wire [31:0] wRegInB23;
wire [31:0] wAIn23;
wire [31:0] wBIn23;
wire [31:0] wRegInA24;
wire [31:0] wRegInB24;
wire [31:0] wAIn24;
wire [31:0] wBIn24;
wire [31:0] wRegInA25;
wire [31:0] wRegInB25;
wire [31:0] wAIn25;
wire [31:0] wBIn25;
wire [31:0] wRegInA26;
wire [31:0] wRegInB26;
wire [31:0] wAIn26;
wire [31:0] wBIn26;
wire [31:0] wRegInA27;
wire [31:0] wRegInB27;
wire [31:0] wAIn27;
wire [31:0] wBIn27;
wire [31:0] wRegInA28;
wire [31:0] wRegInB28;
wire [31:0] wAIn28;
wire [31:0] wBIn28;
wire [31:0] wRegInA29;
wire [31:0] wRegInB29;
wire [31:0] wAIn29;
wire [31:0] wBIn29;
wire [31:0] wRegInA30;
wire [31:0] wRegInB30;
wire [31:0] wAIn30;
wire [31:0] wBIn30;
wire [31:0] wRegInA31;
wire [31:0] wRegInB31;
wire [31:0] wAIn31;
wire [31:0] wBIn31;
wire [31:0] wRegInA32;
wire [31:0] wRegInB32;
wire [31:0] wAIn32;
wire [31:0] wBIn32;
wire [31:0] wRegInA33;
wire [31:0] wRegInB33;
wire [31:0] wAIn33;
wire [31:0] wBIn33;
wire [31:0] wRegInA34;
wire [31:0] wRegInB34;
wire [31:0] wAIn34;
wire [31:0] wBIn34;
wire [31:0] wRegInA35;
wire [31:0] wRegInB35;
wire [31:0] wAIn35;
wire [31:0] wBIn35;
wire [31:0] wRegInA36;
wire [31:0] wRegInB36;
wire [31:0] wAIn36;
wire [31:0] wBIn36;
wire [31:0] wRegInA37;
wire [31:0] wRegInB37;
wire [31:0] wAIn37;
wire [31:0] wBIn37;
wire [31:0] wRegInA38;
wire [31:0] wRegInB38;
wire [31:0] wAIn38;
wire [31:0] wBIn38;
wire [31:0] wRegInA39;
wire [31:0] wRegInB39;
wire [31:0] wAIn39;
wire [31:0] wBIn39;
wire [31:0] wRegInA40;
wire [31:0] wRegInB40;
wire [31:0] wAIn40;
wire [31:0] wBIn40;
wire [31:0] wRegInA41;
wire [31:0] wRegInB41;
wire [31:0] wAIn41;
wire [31:0] wBIn41;
wire [31:0] wRegInA42;
wire [31:0] wRegInB42;
wire [31:0] wAIn42;
wire [31:0] wBIn42;
wire [31:0] wRegInA43;
wire [31:0] wRegInB43;
wire [31:0] wAIn43;
wire [31:0] wBIn43;
wire [31:0] wRegInA44;
wire [31:0] wRegInB44;
wire [31:0] wAIn44;
wire [31:0] wBIn44;
wire [31:0] wRegInA45;
wire [31:0] wRegInB45;
wire [31:0] wAIn45;
wire [31:0] wBIn45;
wire [31:0] wRegInA46;
wire [31:0] wRegInB46;
wire [31:0] wAIn46;
wire [31:0] wBIn46;
wire [31:0] wRegInA47;
wire [31:0] wRegInB47;
wire [31:0] wAIn47;
wire [31:0] wBIn47;
wire [31:0] wRegInA48;
wire [31:0] wRegInB48;
wire [31:0] wAIn48;
wire [31:0] wBIn48;
wire [31:0] wRegInA49;
wire [31:0] wRegInB49;
wire [31:0] wAIn49;
wire [31:0] wBIn49;
wire [31:0] wRegInA50;
wire [31:0] wRegInB50;
wire [31:0] wAIn50;
wire [31:0] wBIn50;
wire [31:0] wRegInA51;
wire [31:0] wRegInB51;
wire [31:0] wAIn51;
wire [31:0] wBIn51;
wire [31:0] wRegInA52;
wire [31:0] wRegInB52;
wire [31:0] wAIn52;
wire [31:0] wBIn52;
wire [31:0] wRegInA53;
wire [31:0] wRegInB53;
wire [31:0] wAIn53;
wire [31:0] wBIn53;
wire [31:0] wRegInA54;
wire [31:0] wRegInB54;
wire [31:0] wAIn54;
wire [31:0] wBIn54;
wire [31:0] wRegInA55;
wire [31:0] wRegInB55;
wire [31:0] wAIn55;
wire [31:0] wBIn55;
wire [31:0] wRegInA56;
wire [31:0] wRegInB56;
wire [31:0] wAIn56;
wire [31:0] wBIn56;
wire [31:0] wRegInA57;
wire [31:0] wRegInB57;
wire [31:0] wAIn57;
wire [31:0] wBIn57;
wire [31:0] wRegInA58;
wire [31:0] wRegInB58;
wire [31:0] wAIn58;
wire [31:0] wBIn58;
wire [31:0] wRegInA59;
wire [31:0] wRegInB59;
wire [31:0] wAIn59;
wire [31:0] wBIn59;
wire [31:0] wRegInA60;
wire [31:0] wRegInB60;
wire [31:0] wAIn60;
wire [31:0] wBIn60;
wire [31:0] wRegInA61;
wire [31:0] wRegInB61;
wire [31:0] wAIn61;
wire [31:0] wBIn61;
wire [31:0] wRegInA62;
wire [31:0] wRegInB62;
wire [31:0] wAIn62;
wire [31:0] wBIn62;
wire [31:0] wRegInA63;
wire [31:0] wRegInB63;
wire [31:0] wAIn63;
wire [31:0] wBIn63;
wire [31:0] wRegInA64;
wire [31:0] wRegInB64;
wire [31:0] wAIn64;
wire [31:0] wBIn64;
wire [31:0] wRegInA65;
wire [31:0] wRegInB65;
wire [31:0] wAIn65;
wire [31:0] wBIn65;
wire [31:0] wRegInA66;
wire [31:0] wRegInB66;
wire [31:0] wAIn66;
wire [31:0] wBIn66;
wire [31:0] wRegInA67;
wire [31:0] wRegInB67;
wire [31:0] wAIn67;
wire [31:0] wBIn67;
wire [31:0] wRegInA68;
wire [31:0] wRegInB68;
wire [31:0] wAIn68;
wire [31:0] wBIn68;
wire [31:0] wRegInA69;
wire [31:0] wRegInB69;
wire [31:0] wAIn69;
wire [31:0] wBIn69;
wire [31:0] wRegInA70;
wire [31:0] wRegInB70;
wire [31:0] wAIn70;
wire [31:0] wBIn70;
wire [31:0] wRegInA71;
wire [31:0] wRegInB71;
wire [31:0] wAIn71;
wire [31:0] wBIn71;
wire [31:0] wRegInA72;
wire [31:0] wRegInB72;
wire [31:0] wAIn72;
wire [31:0] wBIn72;
wire [31:0] wRegInA73;
wire [31:0] wRegInB73;
wire [31:0] wAIn73;
wire [31:0] wBIn73;
wire [31:0] wRegInA74;
wire [31:0] wRegInB74;
wire [31:0] wAIn74;
wire [31:0] wBIn74;
wire [31:0] wRegInA75;
wire [31:0] wRegInB75;
wire [31:0] wAIn75;
wire [31:0] wBIn75;
wire [31:0] wRegInA76;
wire [31:0] wRegInB76;
wire [31:0] wAIn76;
wire [31:0] wBIn76;
wire [31:0] wRegInA77;
wire [31:0] wRegInB77;
wire [31:0] wAIn77;
wire [31:0] wBIn77;
wire [31:0] wRegInA78;
wire [31:0] wRegInB78;
wire [31:0] wAIn78;
wire [31:0] wBIn78;
wire [31:0] wRegInA79;
wire [31:0] wRegInB79;
wire [31:0] wAIn79;
wire [31:0] wBIn79;
wire [31:0] wRegInA80;
wire [31:0] wRegInB80;
wire [31:0] wAIn80;
wire [31:0] wBIn80;
wire [31:0] wRegInA81;
wire [31:0] wRegInB81;
wire [31:0] wAIn81;
wire [31:0] wBIn81;
wire [31:0] wRegInA82;
wire [31:0] wRegInB82;
wire [31:0] wAIn82;
wire [31:0] wBIn82;
wire [31:0] wRegInA83;
wire [31:0] wRegInB83;
wire [31:0] wAIn83;
wire [31:0] wBIn83;
wire [31:0] wRegInA84;
wire [31:0] wRegInB84;
wire [31:0] wAIn84;
wire [31:0] wBIn84;
wire [31:0] wRegInA85;
wire [31:0] wRegInB85;
wire [31:0] wAIn85;
wire [31:0] wBIn85;
wire [31:0] wRegInA86;
wire [31:0] wRegInB86;
wire [31:0] wAIn86;
wire [31:0] wBIn86;
wire [31:0] wRegInA87;
wire [31:0] wRegInB87;
wire [31:0] wAIn87;
wire [31:0] wBIn87;
wire [31:0] wRegInA88;
wire [31:0] wRegInB88;
wire [31:0] wAIn88;
wire [31:0] wBIn88;
wire [31:0] wRegInA89;
wire [31:0] wRegInB89;
wire [31:0] wAIn89;
wire [31:0] wBIn89;
wire [31:0] wRegInA90;
wire [31:0] wRegInB90;
wire [31:0] wAIn90;
wire [31:0] wBIn90;
wire [31:0] wRegInA91;
wire [31:0] wRegInB91;
wire [31:0] wAIn91;
wire [31:0] wBIn91;
wire [31:0] wRegInA92;
wire [31:0] wRegInB92;
wire [31:0] wAIn92;
wire [31:0] wBIn92;
wire [31:0] wRegInA93;
wire [31:0] wRegInB93;
wire [31:0] wAIn93;
wire [31:0] wBIn93;
wire [31:0] wRegInA94;
wire [31:0] wRegInB94;
wire [31:0] wAIn94;
wire [31:0] wBIn94;
wire [31:0] wRegInA95;
wire [31:0] wRegInB95;
wire [31:0] wAIn95;
wire [31:0] wBIn95;
wire [31:0] wRegInA96;
wire [31:0] wRegInB96;
wire [31:0] wAIn96;
wire [31:0] wBIn96;
wire [31:0] wRegInA97;
wire [31:0] wRegInB97;
wire [31:0] wAIn97;
wire [31:0] wBIn97;
wire [31:0] wRegInA98;
wire [31:0] wRegInB98;
wire [31:0] wAIn98;
wire [31:0] wBIn98;
wire [31:0] wRegInA99;
wire [31:0] wRegInB99;
wire [31:0] wAIn99;
wire [31:0] wBIn99;
wire [31:0] wRegInA100;
wire [31:0] wRegInB100;
wire [31:0] wAIn100;
wire [31:0] wBIn100;
wire [31:0] wRegInA101;
wire [31:0] wRegInB101;
wire [31:0] wAIn101;
wire [31:0] wBIn101;
wire [31:0] wRegInA102;
wire [31:0] wRegInB102;
wire [31:0] wAIn102;
wire [31:0] wBIn102;
wire [31:0] wRegInA103;
wire [31:0] wRegInB103;
wire [31:0] wAIn103;
wire [31:0] wBIn103;
wire [31:0] wRegInA104;
wire [31:0] wRegInB104;
wire [31:0] wAIn104;
wire [31:0] wBIn104;
wire [31:0] wRegInA105;
wire [31:0] wRegInB105;
wire [31:0] wAIn105;
wire [31:0] wBIn105;
wire [31:0] wRegInA106;
wire [31:0] wRegInB106;
wire [31:0] wAIn106;
wire [31:0] wBIn106;
wire [31:0] wRegInA107;
wire [31:0] wRegInB107;
wire [31:0] wAIn107;
wire [31:0] wBIn107;
wire [31:0] wRegInA108;
wire [31:0] wRegInB108;
wire [31:0] wAIn108;
wire [31:0] wBIn108;
wire [31:0] wRegInA109;
wire [31:0] wRegInB109;
wire [31:0] wAIn109;
wire [31:0] wBIn109;
wire [31:0] wRegInA110;
wire [31:0] wRegInB110;
wire [31:0] wAIn110;
wire [31:0] wBIn110;
wire [31:0] wRegInA111;
wire [31:0] wRegInB111;
wire [31:0] wAIn111;
wire [31:0] wBIn111;
wire [31:0] wRegInA112;
wire [31:0] wRegInB112;
wire [31:0] wAIn112;
wire [31:0] wBIn112;
wire [31:0] wRegInA113;
wire [31:0] wRegInB113;
wire [31:0] wAIn113;
wire [31:0] wBIn113;
wire [31:0] wRegInA114;
wire [31:0] wRegInB114;
wire [31:0] wAIn114;
wire [31:0] wBIn114;
wire [31:0] wRegInA115;
wire [31:0] wRegInB115;
wire [31:0] wAIn115;
wire [31:0] wBIn115;
wire [31:0] wRegInA116;
wire [31:0] wRegInB116;
wire [31:0] wAIn116;
wire [31:0] wBIn116;
wire [31:0] wRegInA117;
wire [31:0] wRegInB117;
wire [31:0] wAIn117;
wire [31:0] wBIn117;
wire [31:0] wRegInA118;
wire [31:0] wRegInB118;
wire [31:0] wAIn118;
wire [31:0] wBIn118;
wire [31:0] wRegInA119;
wire [31:0] wRegInB119;
wire [31:0] wAIn119;
wire [31:0] wBIn119;
wire [31:0] wRegInA120;
wire [31:0] wRegInB120;
wire [31:0] wAIn120;
wire [31:0] wBIn120;
wire [31:0] wRegInA121;
wire [31:0] wRegInB121;
wire [31:0] wAIn121;
wire [31:0] wBIn121;
wire [31:0] wRegInA122;
wire [31:0] wRegInB122;
wire [31:0] wAIn122;
wire [31:0] wBIn122;
wire [31:0] wRegInA123;
wire [31:0] wRegInB123;
wire [31:0] wAIn123;
wire [31:0] wBIn123;
wire [31:0] wRegInA124;
wire [31:0] wRegInB124;
wire [31:0] wAIn124;
wire [31:0] wBIn124;
wire [31:0] wRegInA125;
wire [31:0] wRegInB125;
wire [31:0] wAIn125;
wire [31:0] wBIn125;
wire [31:0] wRegInA126;
wire [31:0] wRegInB126;
wire [31:0] wAIn126;
wire [31:0] wBIn126;
wire [31:0] wRegInA127;
wire [31:0] wRegInB127;
wire [31:0] wAIn127;
wire [31:0] wBIn127;
wire [31:0] wAMid0;
wire [31:0] wBMid0;
wire [31:0] wAMid1;
wire [31:0] wBMid1;
wire [31:0] wAMid2;
wire [31:0] wBMid2;
wire [31:0] wAMid3;
wire [31:0] wBMid3;
wire [31:0] wAMid4;
wire [31:0] wBMid4;
wire [31:0] wAMid5;
wire [31:0] wBMid5;
wire [31:0] wAMid6;
wire [31:0] wBMid6;
wire [31:0] wAMid7;
wire [31:0] wBMid7;
wire [31:0] wAMid8;
wire [31:0] wBMid8;
wire [31:0] wAMid9;
wire [31:0] wBMid9;
wire [31:0] wAMid10;
wire [31:0] wBMid10;
wire [31:0] wAMid11;
wire [31:0] wBMid11;
wire [31:0] wAMid12;
wire [31:0] wBMid12;
wire [31:0] wAMid13;
wire [31:0] wBMid13;
wire [31:0] wAMid14;
wire [31:0] wBMid14;
wire [31:0] wAMid15;
wire [31:0] wBMid15;
wire [31:0] wAMid16;
wire [31:0] wBMid16;
wire [31:0] wAMid17;
wire [31:0] wBMid17;
wire [31:0] wAMid18;
wire [31:0] wBMid18;
wire [31:0] wAMid19;
wire [31:0] wBMid19;
wire [31:0] wAMid20;
wire [31:0] wBMid20;
wire [31:0] wAMid21;
wire [31:0] wBMid21;
wire [31:0] wAMid22;
wire [31:0] wBMid22;
wire [31:0] wAMid23;
wire [31:0] wBMid23;
wire [31:0] wAMid24;
wire [31:0] wBMid24;
wire [31:0] wAMid25;
wire [31:0] wBMid25;
wire [31:0] wAMid26;
wire [31:0] wBMid26;
wire [31:0] wAMid27;
wire [31:0] wBMid27;
wire [31:0] wAMid28;
wire [31:0] wBMid28;
wire [31:0] wAMid29;
wire [31:0] wBMid29;
wire [31:0] wAMid30;
wire [31:0] wBMid30;
wire [31:0] wAMid31;
wire [31:0] wBMid31;
wire [31:0] wAMid32;
wire [31:0] wBMid32;
wire [31:0] wAMid33;
wire [31:0] wBMid33;
wire [31:0] wAMid34;
wire [31:0] wBMid34;
wire [31:0] wAMid35;
wire [31:0] wBMid35;
wire [31:0] wAMid36;
wire [31:0] wBMid36;
wire [31:0] wAMid37;
wire [31:0] wBMid37;
wire [31:0] wAMid38;
wire [31:0] wBMid38;
wire [31:0] wAMid39;
wire [31:0] wBMid39;
wire [31:0] wAMid40;
wire [31:0] wBMid40;
wire [31:0] wAMid41;
wire [31:0] wBMid41;
wire [31:0] wAMid42;
wire [31:0] wBMid42;
wire [31:0] wAMid43;
wire [31:0] wBMid43;
wire [31:0] wAMid44;
wire [31:0] wBMid44;
wire [31:0] wAMid45;
wire [31:0] wBMid45;
wire [31:0] wAMid46;
wire [31:0] wBMid46;
wire [31:0] wAMid47;
wire [31:0] wBMid47;
wire [31:0] wAMid48;
wire [31:0] wBMid48;
wire [31:0] wAMid49;
wire [31:0] wBMid49;
wire [31:0] wAMid50;
wire [31:0] wBMid50;
wire [31:0] wAMid51;
wire [31:0] wBMid51;
wire [31:0] wAMid52;
wire [31:0] wBMid52;
wire [31:0] wAMid53;
wire [31:0] wBMid53;
wire [31:0] wAMid54;
wire [31:0] wBMid54;
wire [31:0] wAMid55;
wire [31:0] wBMid55;
wire [31:0] wAMid56;
wire [31:0] wBMid56;
wire [31:0] wAMid57;
wire [31:0] wBMid57;
wire [31:0] wAMid58;
wire [31:0] wBMid58;
wire [31:0] wAMid59;
wire [31:0] wBMid59;
wire [31:0] wAMid60;
wire [31:0] wBMid60;
wire [31:0] wAMid61;
wire [31:0] wBMid61;
wire [31:0] wAMid62;
wire [31:0] wBMid62;
wire [31:0] wAMid63;
wire [31:0] wBMid63;
wire [31:0] wAMid64;
wire [31:0] wBMid64;
wire [31:0] wAMid65;
wire [31:0] wBMid65;
wire [31:0] wAMid66;
wire [31:0] wBMid66;
wire [31:0] wAMid67;
wire [31:0] wBMid67;
wire [31:0] wAMid68;
wire [31:0] wBMid68;
wire [31:0] wAMid69;
wire [31:0] wBMid69;
wire [31:0] wAMid70;
wire [31:0] wBMid70;
wire [31:0] wAMid71;
wire [31:0] wBMid71;
wire [31:0] wAMid72;
wire [31:0] wBMid72;
wire [31:0] wAMid73;
wire [31:0] wBMid73;
wire [31:0] wAMid74;
wire [31:0] wBMid74;
wire [31:0] wAMid75;
wire [31:0] wBMid75;
wire [31:0] wAMid76;
wire [31:0] wBMid76;
wire [31:0] wAMid77;
wire [31:0] wBMid77;
wire [31:0] wAMid78;
wire [31:0] wBMid78;
wire [31:0] wAMid79;
wire [31:0] wBMid79;
wire [31:0] wAMid80;
wire [31:0] wBMid80;
wire [31:0] wAMid81;
wire [31:0] wBMid81;
wire [31:0] wAMid82;
wire [31:0] wBMid82;
wire [31:0] wAMid83;
wire [31:0] wBMid83;
wire [31:0] wAMid84;
wire [31:0] wBMid84;
wire [31:0] wAMid85;
wire [31:0] wBMid85;
wire [31:0] wAMid86;
wire [31:0] wBMid86;
wire [31:0] wAMid87;
wire [31:0] wBMid87;
wire [31:0] wAMid88;
wire [31:0] wBMid88;
wire [31:0] wAMid89;
wire [31:0] wBMid89;
wire [31:0] wAMid90;
wire [31:0] wBMid90;
wire [31:0] wAMid91;
wire [31:0] wBMid91;
wire [31:0] wAMid92;
wire [31:0] wBMid92;
wire [31:0] wAMid93;
wire [31:0] wBMid93;
wire [31:0] wAMid94;
wire [31:0] wBMid94;
wire [31:0] wAMid95;
wire [31:0] wBMid95;
wire [31:0] wAMid96;
wire [31:0] wBMid96;
wire [31:0] wAMid97;
wire [31:0] wBMid97;
wire [31:0] wAMid98;
wire [31:0] wBMid98;
wire [31:0] wAMid99;
wire [31:0] wBMid99;
wire [31:0] wAMid100;
wire [31:0] wBMid100;
wire [31:0] wAMid101;
wire [31:0] wBMid101;
wire [31:0] wAMid102;
wire [31:0] wBMid102;
wire [31:0] wAMid103;
wire [31:0] wBMid103;
wire [31:0] wAMid104;
wire [31:0] wBMid104;
wire [31:0] wAMid105;
wire [31:0] wBMid105;
wire [31:0] wAMid106;
wire [31:0] wBMid106;
wire [31:0] wAMid107;
wire [31:0] wBMid107;
wire [31:0] wAMid108;
wire [31:0] wBMid108;
wire [31:0] wAMid109;
wire [31:0] wBMid109;
wire [31:0] wAMid110;
wire [31:0] wBMid110;
wire [31:0] wAMid111;
wire [31:0] wBMid111;
wire [31:0] wAMid112;
wire [31:0] wBMid112;
wire [31:0] wAMid113;
wire [31:0] wBMid113;
wire [31:0] wAMid114;
wire [31:0] wBMid114;
wire [31:0] wAMid115;
wire [31:0] wBMid115;
wire [31:0] wAMid116;
wire [31:0] wBMid116;
wire [31:0] wAMid117;
wire [31:0] wBMid117;
wire [31:0] wAMid118;
wire [31:0] wBMid118;
wire [31:0] wAMid119;
wire [31:0] wBMid119;
wire [31:0] wAMid120;
wire [31:0] wBMid120;
wire [31:0] wAMid121;
wire [31:0] wBMid121;
wire [31:0] wAMid122;
wire [31:0] wBMid122;
wire [31:0] wAMid123;
wire [31:0] wBMid123;
wire [31:0] wAMid124;
wire [31:0] wBMid124;
wire [31:0] wAMid125;
wire [31:0] wBMid125;
wire [31:0] wAMid126;
wire [31:0] wBMid126;
wire [0:0] wEnable;
wire [0:0] ScanEnable;
wire [31:0] ScanLink0;
wire [31:0] ScanLink1;
wire [31:0] ScanLink2;
wire [31:0] ScanLink3;
wire [31:0] ScanLink4;
wire [31:0] ScanLink5;
wire [31:0] ScanLink6;
wire [31:0] ScanLink7;
wire [31:0] ScanLink8;
wire [31:0] ScanLink9;
wire [31:0] ScanLink10;
wire [31:0] ScanLink11;
wire [31:0] ScanLink12;
wire [31:0] ScanLink13;
wire [31:0] ScanLink14;
wire [31:0] ScanLink15;
wire [31:0] ScanLink16;
wire [31:0] ScanLink17;
wire [31:0] ScanLink18;
wire [31:0] ScanLink19;
wire [31:0] ScanLink20;
wire [31:0] ScanLink21;
wire [31:0] ScanLink22;
wire [31:0] ScanLink23;
wire [31:0] ScanLink24;
wire [31:0] ScanLink25;
wire [31:0] ScanLink26;
wire [31:0] ScanLink27;
wire [31:0] ScanLink28;
wire [31:0] ScanLink29;
wire [31:0] ScanLink30;
wire [31:0] ScanLink31;
wire [31:0] ScanLink32;
wire [31:0] ScanLink33;
wire [31:0] ScanLink34;
wire [31:0] ScanLink35;
wire [31:0] ScanLink36;
wire [31:0] ScanLink37;
wire [31:0] ScanLink38;
wire [31:0] ScanLink39;
wire [31:0] ScanLink40;
wire [31:0] ScanLink41;
wire [31:0] ScanLink42;
wire [31:0] ScanLink43;
wire [31:0] ScanLink44;
wire [31:0] ScanLink45;
wire [31:0] ScanLink46;
wire [31:0] ScanLink47;
wire [31:0] ScanLink48;
wire [31:0] ScanLink49;
wire [31:0] ScanLink50;
wire [31:0] ScanLink51;
wire [31:0] ScanLink52;
wire [31:0] ScanLink53;
wire [31:0] ScanLink54;
wire [31:0] ScanLink55;
wire [31:0] ScanLink56;
wire [31:0] ScanLink57;
wire [31:0] ScanLink58;
wire [31:0] ScanLink59;
wire [31:0] ScanLink60;
wire [31:0] ScanLink61;
wire [31:0] ScanLink62;
wire [31:0] ScanLink63;
wire [31:0] ScanLink64;
wire [31:0] ScanLink65;
wire [31:0] ScanLink66;
wire [31:0] ScanLink67;
wire [31:0] ScanLink68;
wire [31:0] ScanLink69;
wire [31:0] ScanLink70;
wire [31:0] ScanLink71;
wire [31:0] ScanLink72;
wire [31:0] ScanLink73;
wire [31:0] ScanLink74;
wire [31:0] ScanLink75;
wire [31:0] ScanLink76;
wire [31:0] ScanLink77;
wire [31:0] ScanLink78;
wire [31:0] ScanLink79;
wire [31:0] ScanLink80;
wire [31:0] ScanLink81;
wire [31:0] ScanLink82;
wire [31:0] ScanLink83;
wire [31:0] ScanLink84;
wire [31:0] ScanLink85;
wire [31:0] ScanLink86;
wire [31:0] ScanLink87;
wire [31:0] ScanLink88;
wire [31:0] ScanLink89;
wire [31:0] ScanLink90;
wire [31:0] ScanLink91;
wire [31:0] ScanLink92;
wire [31:0] ScanLink93;
wire [31:0] ScanLink94;
wire [31:0] ScanLink95;
wire [31:0] ScanLink96;
wire [31:0] ScanLink97;
wire [31:0] ScanLink98;
wire [31:0] ScanLink99;
wire [31:0] ScanLink100;
wire [31:0] ScanLink101;
wire [31:0] ScanLink102;
wire [31:0] ScanLink103;
wire [31:0] ScanLink104;
wire [31:0] ScanLink105;
wire [31:0] ScanLink106;
wire [31:0] ScanLink107;
wire [31:0] ScanLink108;
wire [31:0] ScanLink109;
wire [31:0] ScanLink110;
wire [31:0] ScanLink111;
wire [31:0] ScanLink112;
wire [31:0] ScanLink113;
wire [31:0] ScanLink114;
wire [31:0] ScanLink115;
wire [31:0] ScanLink116;
wire [31:0] ScanLink117;
wire [31:0] ScanLink118;
wire [31:0] ScanLink119;
wire [31:0] ScanLink120;
wire [31:0] ScanLink121;
wire [31:0] ScanLink122;
wire [31:0] ScanLink123;
wire [31:0] ScanLink124;
wire [31:0] ScanLink125;
wire [31:0] ScanLink126;
wire [31:0] ScanLink127;
wire [31:0] ScanLink128;
wire [31:0] ScanLink129;
wire [31:0] ScanLink130;
wire [31:0] ScanLink131;
wire [31:0] ScanLink132;
wire [31:0] ScanLink133;
wire [31:0] ScanLink134;
wire [31:0] ScanLink135;
wire [31:0] ScanLink136;
wire [31:0] ScanLink137;
wire [31:0] ScanLink138;
wire [31:0] ScanLink139;
wire [31:0] ScanLink140;
wire [31:0] ScanLink141;
wire [31:0] ScanLink142;
wire [31:0] ScanLink143;
wire [31:0] ScanLink144;
wire [31:0] ScanLink145;
wire [31:0] ScanLink146;
wire [31:0] ScanLink147;
wire [31:0] ScanLink148;
wire [31:0] ScanLink149;
wire [31:0] ScanLink150;
wire [31:0] ScanLink151;
wire [31:0] ScanLink152;
wire [31:0] ScanLink153;
wire [31:0] ScanLink154;
wire [31:0] ScanLink155;
wire [31:0] ScanLink156;
wire [31:0] ScanLink157;
wire [31:0] ScanLink158;
wire [31:0] ScanLink159;
wire [31:0] ScanLink160;
wire [31:0] ScanLink161;
wire [31:0] ScanLink162;
wire [31:0] ScanLink163;
wire [31:0] ScanLink164;
wire [31:0] ScanLink165;
wire [31:0] ScanLink166;
wire [31:0] ScanLink167;
wire [31:0] ScanLink168;
wire [31:0] ScanLink169;
wire [31:0] ScanLink170;
wire [31:0] ScanLink171;
wire [31:0] ScanLink172;
wire [31:0] ScanLink173;
wire [31:0] ScanLink174;
wire [31:0] ScanLink175;
wire [31:0] ScanLink176;
wire [31:0] ScanLink177;
wire [31:0] ScanLink178;
wire [31:0] ScanLink179;
wire [31:0] ScanLink180;
wire [31:0] ScanLink181;
wire [31:0] ScanLink182;
wire [31:0] ScanLink183;
wire [31:0] ScanLink184;
wire [31:0] ScanLink185;
wire [31:0] ScanLink186;
wire [31:0] ScanLink187;
wire [31:0] ScanLink188;
wire [31:0] ScanLink189;
wire [31:0] ScanLink190;
wire [31:0] ScanLink191;
wire [31:0] ScanLink192;
wire [31:0] ScanLink193;
wire [31:0] ScanLink194;
wire [31:0] ScanLink195;
wire [31:0] ScanLink196;
wire [31:0] ScanLink197;
wire [31:0] ScanLink198;
wire [31:0] ScanLink199;
wire [31:0] ScanLink200;
wire [31:0] ScanLink201;
wire [31:0] ScanLink202;
wire [31:0] ScanLink203;
wire [31:0] ScanLink204;
wire [31:0] ScanLink205;
wire [31:0] ScanLink206;
wire [31:0] ScanLink207;
wire [31:0] ScanLink208;
wire [31:0] ScanLink209;
wire [31:0] ScanLink210;
wire [31:0] ScanLink211;
wire [31:0] ScanLink212;
wire [31:0] ScanLink213;
wire [31:0] ScanLink214;
wire [31:0] ScanLink215;
wire [31:0] ScanLink216;
wire [31:0] ScanLink217;
wire [31:0] ScanLink218;
wire [31:0] ScanLink219;
wire [31:0] ScanLink220;
wire [31:0] ScanLink221;
wire [31:0] ScanLink222;
wire [31:0] ScanLink223;
wire [31:0] ScanLink224;
wire [31:0] ScanLink225;
wire [31:0] ScanLink226;
wire [31:0] ScanLink227;
wire [31:0] ScanLink228;
wire [31:0] ScanLink229;
wire [31:0] ScanLink230;
wire [31:0] ScanLink231;
wire [31:0] ScanLink232;
wire [31:0] ScanLink233;
wire [31:0] ScanLink234;
wire [31:0] ScanLink235;
wire [31:0] ScanLink236;
wire [31:0] ScanLink237;
wire [31:0] ScanLink238;
wire [31:0] ScanLink239;
wire [31:0] ScanLink240;
wire [31:0] ScanLink241;
wire [31:0] ScanLink242;
wire [31:0] ScanLink243;
wire [31:0] ScanLink244;
wire [31:0] ScanLink245;
wire [31:0] ScanLink246;
wire [31:0] ScanLink247;
wire [31:0] ScanLink248;
wire [31:0] ScanLink249;
wire [31:0] ScanLink250;
wire [31:0] ScanLink251;
wire [31:0] ScanLink252;
wire [31:0] ScanLink253;
wire [31:0] ScanLink254;
wire [31:0] ScanLink255;
wire [31:0] ScanLink256;
BubbleSort_Node #( 32 ) BSN1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn0), .BIn(wBIn0), .HiOut(wRegInA0), .LoOut(wAMid0) );
BubbleSort_Node #( 32 ) BSN1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn1), .BIn(wBIn1), .HiOut(wBMid0), .LoOut(wAMid1) );
BubbleSort_Node #( 32 ) BSN1_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn2), .BIn(wBIn2), .HiOut(wBMid1), .LoOut(wAMid2) );
BubbleSort_Node #( 32 ) BSN1_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn3), .BIn(wBIn3), .HiOut(wBMid2), .LoOut(wAMid3) );
BubbleSort_Node #( 32 ) BSN1_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn4), .BIn(wBIn4), .HiOut(wBMid3), .LoOut(wAMid4) );
BubbleSort_Node #( 32 ) BSN1_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn5), .BIn(wBIn5), .HiOut(wBMid4), .LoOut(wAMid5) );
BubbleSort_Node #( 32 ) BSN1_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn6), .BIn(wBIn6), .HiOut(wBMid5), .LoOut(wAMid6) );
BubbleSort_Node #( 32 ) BSN1_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn7), .BIn(wBIn7), .HiOut(wBMid6), .LoOut(wAMid7) );
BubbleSort_Node #( 32 ) BSN1_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn8), .BIn(wBIn8), .HiOut(wBMid7), .LoOut(wAMid8) );
BubbleSort_Node #( 32 ) BSN1_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn9), .BIn(wBIn9), .HiOut(wBMid8), .LoOut(wAMid9) );
BubbleSort_Node #( 32 ) BSN1_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn10), .BIn(wBIn10), .HiOut(wBMid9), .LoOut(wAMid10) );
BubbleSort_Node #( 32 ) BSN1_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn11), .BIn(wBIn11), .HiOut(wBMid10), .LoOut(wAMid11) );
BubbleSort_Node #( 32 ) BSN1_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn12), .BIn(wBIn12), .HiOut(wBMid11), .LoOut(wAMid12) );
BubbleSort_Node #( 32 ) BSN1_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn13), .BIn(wBIn13), .HiOut(wBMid12), .LoOut(wAMid13) );
BubbleSort_Node #( 32 ) BSN1_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn14), .BIn(wBIn14), .HiOut(wBMid13), .LoOut(wAMid14) );
BubbleSort_Node #( 32 ) BSN1_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn15), .BIn(wBIn15), .HiOut(wBMid14), .LoOut(wAMid15) );
BubbleSort_Node #( 32 ) BSN1_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn16), .BIn(wBIn16), .HiOut(wBMid15), .LoOut(wAMid16) );
BubbleSort_Node #( 32 ) BSN1_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn17), .BIn(wBIn17), .HiOut(wBMid16), .LoOut(wAMid17) );
BubbleSort_Node #( 32 ) BSN1_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn18), .BIn(wBIn18), .HiOut(wBMid17), .LoOut(wAMid18) );
BubbleSort_Node #( 32 ) BSN1_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn19), .BIn(wBIn19), .HiOut(wBMid18), .LoOut(wAMid19) );
BubbleSort_Node #( 32 ) BSN1_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn20), .BIn(wBIn20), .HiOut(wBMid19), .LoOut(wAMid20) );
BubbleSort_Node #( 32 ) BSN1_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn21), .BIn(wBIn21), .HiOut(wBMid20), .LoOut(wAMid21) );
BubbleSort_Node #( 32 ) BSN1_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn22), .BIn(wBIn22), .HiOut(wBMid21), .LoOut(wAMid22) );
BubbleSort_Node #( 32 ) BSN1_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn23), .BIn(wBIn23), .HiOut(wBMid22), .LoOut(wAMid23) );
BubbleSort_Node #( 32 ) BSN1_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn24), .BIn(wBIn24), .HiOut(wBMid23), .LoOut(wAMid24) );
BubbleSort_Node #( 32 ) BSN1_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn25), .BIn(wBIn25), .HiOut(wBMid24), .LoOut(wAMid25) );
BubbleSort_Node #( 32 ) BSN1_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn26), .BIn(wBIn26), .HiOut(wBMid25), .LoOut(wAMid26) );
BubbleSort_Node #( 32 ) BSN1_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn27), .BIn(wBIn27), .HiOut(wBMid26), .LoOut(wAMid27) );
BubbleSort_Node #( 32 ) BSN1_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn28), .BIn(wBIn28), .HiOut(wBMid27), .LoOut(wAMid28) );
BubbleSort_Node #( 32 ) BSN1_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn29), .BIn(wBIn29), .HiOut(wBMid28), .LoOut(wAMid29) );
BubbleSort_Node #( 32 ) BSN1_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn30), .BIn(wBIn30), .HiOut(wBMid29), .LoOut(wAMid30) );
BubbleSort_Node #( 32 ) BSN1_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn31), .BIn(wBIn31), .HiOut(wBMid30), .LoOut(wAMid31) );
BubbleSort_Node #( 32 ) BSN1_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn32), .BIn(wBIn32), .HiOut(wBMid31), .LoOut(wAMid32) );
BubbleSort_Node #( 32 ) BSN1_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn33), .BIn(wBIn33), .HiOut(wBMid32), .LoOut(wAMid33) );
BubbleSort_Node #( 32 ) BSN1_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn34), .BIn(wBIn34), .HiOut(wBMid33), .LoOut(wAMid34) );
BubbleSort_Node #( 32 ) BSN1_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn35), .BIn(wBIn35), .HiOut(wBMid34), .LoOut(wAMid35) );
BubbleSort_Node #( 32 ) BSN1_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn36), .BIn(wBIn36), .HiOut(wBMid35), .LoOut(wAMid36) );
BubbleSort_Node #( 32 ) BSN1_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn37), .BIn(wBIn37), .HiOut(wBMid36), .LoOut(wAMid37) );
BubbleSort_Node #( 32 ) BSN1_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn38), .BIn(wBIn38), .HiOut(wBMid37), .LoOut(wAMid38) );
BubbleSort_Node #( 32 ) BSN1_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn39), .BIn(wBIn39), .HiOut(wBMid38), .LoOut(wAMid39) );
BubbleSort_Node #( 32 ) BSN1_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn40), .BIn(wBIn40), .HiOut(wBMid39), .LoOut(wAMid40) );
BubbleSort_Node #( 32 ) BSN1_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn41), .BIn(wBIn41), .HiOut(wBMid40), .LoOut(wAMid41) );
BubbleSort_Node #( 32 ) BSN1_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn42), .BIn(wBIn42), .HiOut(wBMid41), .LoOut(wAMid42) );
BubbleSort_Node #( 32 ) BSN1_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn43), .BIn(wBIn43), .HiOut(wBMid42), .LoOut(wAMid43) );
BubbleSort_Node #( 32 ) BSN1_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn44), .BIn(wBIn44), .HiOut(wBMid43), .LoOut(wAMid44) );
BubbleSort_Node #( 32 ) BSN1_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn45), .BIn(wBIn45), .HiOut(wBMid44), .LoOut(wAMid45) );
BubbleSort_Node #( 32 ) BSN1_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn46), .BIn(wBIn46), .HiOut(wBMid45), .LoOut(wAMid46) );
BubbleSort_Node #( 32 ) BSN1_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn47), .BIn(wBIn47), .HiOut(wBMid46), .LoOut(wAMid47) );
BubbleSort_Node #( 32 ) BSN1_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn48), .BIn(wBIn48), .HiOut(wBMid47), .LoOut(wAMid48) );
BubbleSort_Node #( 32 ) BSN1_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn49), .BIn(wBIn49), .HiOut(wBMid48), .LoOut(wAMid49) );
BubbleSort_Node #( 32 ) BSN1_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn50), .BIn(wBIn50), .HiOut(wBMid49), .LoOut(wAMid50) );
BubbleSort_Node #( 32 ) BSN1_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn51), .BIn(wBIn51), .HiOut(wBMid50), .LoOut(wAMid51) );
BubbleSort_Node #( 32 ) BSN1_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn52), .BIn(wBIn52), .HiOut(wBMid51), .LoOut(wAMid52) );
BubbleSort_Node #( 32 ) BSN1_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn53), .BIn(wBIn53), .HiOut(wBMid52), .LoOut(wAMid53) );
BubbleSort_Node #( 32 ) BSN1_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn54), .BIn(wBIn54), .HiOut(wBMid53), .LoOut(wAMid54) );
BubbleSort_Node #( 32 ) BSN1_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn55), .BIn(wBIn55), .HiOut(wBMid54), .LoOut(wAMid55) );
BubbleSort_Node #( 32 ) BSN1_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn56), .BIn(wBIn56), .HiOut(wBMid55), .LoOut(wAMid56) );
BubbleSort_Node #( 32 ) BSN1_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn57), .BIn(wBIn57), .HiOut(wBMid56), .LoOut(wAMid57) );
BubbleSort_Node #( 32 ) BSN1_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn58), .BIn(wBIn58), .HiOut(wBMid57), .LoOut(wAMid58) );
BubbleSort_Node #( 32 ) BSN1_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn59), .BIn(wBIn59), .HiOut(wBMid58), .LoOut(wAMid59) );
BubbleSort_Node #( 32 ) BSN1_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn60), .BIn(wBIn60), .HiOut(wBMid59), .LoOut(wAMid60) );
BubbleSort_Node #( 32 ) BSN1_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn61), .BIn(wBIn61), .HiOut(wBMid60), .LoOut(wAMid61) );
BubbleSort_Node #( 32 ) BSN1_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn62), .BIn(wBIn62), .HiOut(wBMid61), .LoOut(wAMid62) );
BubbleSort_Node #( 32 ) BSN1_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn63), .BIn(wBIn63), .HiOut(wBMid62), .LoOut(wAMid63) );
BubbleSort_Node #( 32 ) BSN1_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn64), .BIn(wBIn64), .HiOut(wBMid63), .LoOut(wAMid64) );
BubbleSort_Node #( 32 ) BSN1_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn65), .BIn(wBIn65), .HiOut(wBMid64), .LoOut(wAMid65) );
BubbleSort_Node #( 32 ) BSN1_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn66), .BIn(wBIn66), .HiOut(wBMid65), .LoOut(wAMid66) );
BubbleSort_Node #( 32 ) BSN1_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn67), .BIn(wBIn67), .HiOut(wBMid66), .LoOut(wAMid67) );
BubbleSort_Node #( 32 ) BSN1_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn68), .BIn(wBIn68), .HiOut(wBMid67), .LoOut(wAMid68) );
BubbleSort_Node #( 32 ) BSN1_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn69), .BIn(wBIn69), .HiOut(wBMid68), .LoOut(wAMid69) );
BubbleSort_Node #( 32 ) BSN1_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn70), .BIn(wBIn70), .HiOut(wBMid69), .LoOut(wAMid70) );
BubbleSort_Node #( 32 ) BSN1_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn71), .BIn(wBIn71), .HiOut(wBMid70), .LoOut(wAMid71) );
BubbleSort_Node #( 32 ) BSN1_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn72), .BIn(wBIn72), .HiOut(wBMid71), .LoOut(wAMid72) );
BubbleSort_Node #( 32 ) BSN1_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn73), .BIn(wBIn73), .HiOut(wBMid72), .LoOut(wAMid73) );
BubbleSort_Node #( 32 ) BSN1_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn74), .BIn(wBIn74), .HiOut(wBMid73), .LoOut(wAMid74) );
BubbleSort_Node #( 32 ) BSN1_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn75), .BIn(wBIn75), .HiOut(wBMid74), .LoOut(wAMid75) );
BubbleSort_Node #( 32 ) BSN1_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn76), .BIn(wBIn76), .HiOut(wBMid75), .LoOut(wAMid76) );
BubbleSort_Node #( 32 ) BSN1_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn77), .BIn(wBIn77), .HiOut(wBMid76), .LoOut(wAMid77) );
BubbleSort_Node #( 32 ) BSN1_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn78), .BIn(wBIn78), .HiOut(wBMid77), .LoOut(wAMid78) );
BubbleSort_Node #( 32 ) BSN1_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn79), .BIn(wBIn79), .HiOut(wBMid78), .LoOut(wAMid79) );
BubbleSort_Node #( 32 ) BSN1_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn80), .BIn(wBIn80), .HiOut(wBMid79), .LoOut(wAMid80) );
BubbleSort_Node #( 32 ) BSN1_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn81), .BIn(wBIn81), .HiOut(wBMid80), .LoOut(wAMid81) );
BubbleSort_Node #( 32 ) BSN1_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn82), .BIn(wBIn82), .HiOut(wBMid81), .LoOut(wAMid82) );
BubbleSort_Node #( 32 ) BSN1_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn83), .BIn(wBIn83), .HiOut(wBMid82), .LoOut(wAMid83) );
BubbleSort_Node #( 32 ) BSN1_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn84), .BIn(wBIn84), .HiOut(wBMid83), .LoOut(wAMid84) );
BubbleSort_Node #( 32 ) BSN1_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn85), .BIn(wBIn85), .HiOut(wBMid84), .LoOut(wAMid85) );
BubbleSort_Node #( 32 ) BSN1_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn86), .BIn(wBIn86), .HiOut(wBMid85), .LoOut(wAMid86) );
BubbleSort_Node #( 32 ) BSN1_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn87), .BIn(wBIn87), .HiOut(wBMid86), .LoOut(wAMid87) );
BubbleSort_Node #( 32 ) BSN1_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn88), .BIn(wBIn88), .HiOut(wBMid87), .LoOut(wAMid88) );
BubbleSort_Node #( 32 ) BSN1_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn89), .BIn(wBIn89), .HiOut(wBMid88), .LoOut(wAMid89) );
BubbleSort_Node #( 32 ) BSN1_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn90), .BIn(wBIn90), .HiOut(wBMid89), .LoOut(wAMid90) );
BubbleSort_Node #( 32 ) BSN1_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn91), .BIn(wBIn91), .HiOut(wBMid90), .LoOut(wAMid91) );
BubbleSort_Node #( 32 ) BSN1_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn92), .BIn(wBIn92), .HiOut(wBMid91), .LoOut(wAMid92) );
BubbleSort_Node #( 32 ) BSN1_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn93), .BIn(wBIn93), .HiOut(wBMid92), .LoOut(wAMid93) );
BubbleSort_Node #( 32 ) BSN1_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn94), .BIn(wBIn94), .HiOut(wBMid93), .LoOut(wAMid94) );
BubbleSort_Node #( 32 ) BSN1_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn95), .BIn(wBIn95), .HiOut(wBMid94), .LoOut(wAMid95) );
BubbleSort_Node #( 32 ) BSN1_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn96), .BIn(wBIn96), .HiOut(wBMid95), .LoOut(wAMid96) );
BubbleSort_Node #( 32 ) BSN1_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn97), .BIn(wBIn97), .HiOut(wBMid96), .LoOut(wAMid97) );
BubbleSort_Node #( 32 ) BSN1_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn98), .BIn(wBIn98), .HiOut(wBMid97), .LoOut(wAMid98) );
BubbleSort_Node #( 32 ) BSN1_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn99), .BIn(wBIn99), .HiOut(wBMid98), .LoOut(wAMid99) );
BubbleSort_Node #( 32 ) BSN1_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn100), .BIn(wBIn100), .HiOut(wBMid99), .LoOut(wAMid100) );
BubbleSort_Node #( 32 ) BSN1_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn101), .BIn(wBIn101), .HiOut(wBMid100), .LoOut(wAMid101) );
BubbleSort_Node #( 32 ) BSN1_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn102), .BIn(wBIn102), .HiOut(wBMid101), .LoOut(wAMid102) );
BubbleSort_Node #( 32 ) BSN1_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn103), .BIn(wBIn103), .HiOut(wBMid102), .LoOut(wAMid103) );
BubbleSort_Node #( 32 ) BSN1_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn104), .BIn(wBIn104), .HiOut(wBMid103), .LoOut(wAMid104) );
BubbleSort_Node #( 32 ) BSN1_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn105), .BIn(wBIn105), .HiOut(wBMid104), .LoOut(wAMid105) );
BubbleSort_Node #( 32 ) BSN1_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn106), .BIn(wBIn106), .HiOut(wBMid105), .LoOut(wAMid106) );
BubbleSort_Node #( 32 ) BSN1_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn107), .BIn(wBIn107), .HiOut(wBMid106), .LoOut(wAMid107) );
BubbleSort_Node #( 32 ) BSN1_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn108), .BIn(wBIn108), .HiOut(wBMid107), .LoOut(wAMid108) );
BubbleSort_Node #( 32 ) BSN1_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn109), .BIn(wBIn109), .HiOut(wBMid108), .LoOut(wAMid109) );
BubbleSort_Node #( 32 ) BSN1_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn110), .BIn(wBIn110), .HiOut(wBMid109), .LoOut(wAMid110) );
BubbleSort_Node #( 32 ) BSN1_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn111), .BIn(wBIn111), .HiOut(wBMid110), .LoOut(wAMid111) );
BubbleSort_Node #( 32 ) BSN1_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn112), .BIn(wBIn112), .HiOut(wBMid111), .LoOut(wAMid112) );
BubbleSort_Node #( 32 ) BSN1_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn113), .BIn(wBIn113), .HiOut(wBMid112), .LoOut(wAMid113) );
BubbleSort_Node #( 32 ) BSN1_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn114), .BIn(wBIn114), .HiOut(wBMid113), .LoOut(wAMid114) );
BubbleSort_Node #( 32 ) BSN1_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn115), .BIn(wBIn115), .HiOut(wBMid114), .LoOut(wAMid115) );
BubbleSort_Node #( 32 ) BSN1_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn116), .BIn(wBIn116), .HiOut(wBMid115), .LoOut(wAMid116) );
BubbleSort_Node #( 32 ) BSN1_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn117), .BIn(wBIn117), .HiOut(wBMid116), .LoOut(wAMid117) );
BubbleSort_Node #( 32 ) BSN1_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn118), .BIn(wBIn118), .HiOut(wBMid117), .LoOut(wAMid118) );
BubbleSort_Node #( 32 ) BSN1_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn119), .BIn(wBIn119), .HiOut(wBMid118), .LoOut(wAMid119) );
BubbleSort_Node #( 32 ) BSN1_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn120), .BIn(wBIn120), .HiOut(wBMid119), .LoOut(wAMid120) );
BubbleSort_Node #( 32 ) BSN1_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn121), .BIn(wBIn121), .HiOut(wBMid120), .LoOut(wAMid121) );
BubbleSort_Node #( 32 ) BSN1_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn122), .BIn(wBIn122), .HiOut(wBMid121), .LoOut(wAMid122) );
BubbleSort_Node #( 32 ) BSN1_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn123), .BIn(wBIn123), .HiOut(wBMid122), .LoOut(wAMid123) );
BubbleSort_Node #( 32 ) BSN1_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn124), .BIn(wBIn124), .HiOut(wBMid123), .LoOut(wAMid124) );
BubbleSort_Node #( 32 ) BSN1_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn125), .BIn(wBIn125), .HiOut(wBMid124), .LoOut(wAMid125) );
BubbleSort_Node #( 32 ) BSN1_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn126), .BIn(wBIn126), .HiOut(wBMid125), .LoOut(wAMid126) );
BubbleSort_Node #( 32 ) BSN1_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn127), .BIn(wBIn127), .HiOut(wBMid126), .LoOut(wRegInB127) );
BubbleSort_Node #( 32 ) BSN2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid0), .BIn(wBMid0), .HiOut(wRegInB0), .LoOut(wRegInA1) );
BubbleSort_Node #( 32 ) BSN2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid1), .BIn(wBMid1), .HiOut(wRegInB1), .LoOut(wRegInA2) );
BubbleSort_Node #( 32 ) BSN2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid2), .BIn(wBMid2), .HiOut(wRegInB2), .LoOut(wRegInA3) );
BubbleSort_Node #( 32 ) BSN2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid3), .BIn(wBMid3), .HiOut(wRegInB3), .LoOut(wRegInA4) );
BubbleSort_Node #( 32 ) BSN2_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid4), .BIn(wBMid4), .HiOut(wRegInB4), .LoOut(wRegInA5) );
BubbleSort_Node #( 32 ) BSN2_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid5), .BIn(wBMid5), .HiOut(wRegInB5), .LoOut(wRegInA6) );
BubbleSort_Node #( 32 ) BSN2_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid6), .BIn(wBMid6), .HiOut(wRegInB6), .LoOut(wRegInA7) );
BubbleSort_Node #( 32 ) BSN2_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid7), .BIn(wBMid7), .HiOut(wRegInB7), .LoOut(wRegInA8) );
BubbleSort_Node #( 32 ) BSN2_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid8), .BIn(wBMid8), .HiOut(wRegInB8), .LoOut(wRegInA9) );
BubbleSort_Node #( 32 ) BSN2_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid9), .BIn(wBMid9), .HiOut(wRegInB9), .LoOut(wRegInA10) );
BubbleSort_Node #( 32 ) BSN2_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid10), .BIn(wBMid10), .HiOut(wRegInB10), .LoOut(wRegInA11) );
BubbleSort_Node #( 32 ) BSN2_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid11), .BIn(wBMid11), .HiOut(wRegInB11), .LoOut(wRegInA12) );
BubbleSort_Node #( 32 ) BSN2_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid12), .BIn(wBMid12), .HiOut(wRegInB12), .LoOut(wRegInA13) );
BubbleSort_Node #( 32 ) BSN2_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid13), .BIn(wBMid13), .HiOut(wRegInB13), .LoOut(wRegInA14) );
BubbleSort_Node #( 32 ) BSN2_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid14), .BIn(wBMid14), .HiOut(wRegInB14), .LoOut(wRegInA15) );
BubbleSort_Node #( 32 ) BSN2_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid15), .BIn(wBMid15), .HiOut(wRegInB15), .LoOut(wRegInA16) );
BubbleSort_Node #( 32 ) BSN2_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid16), .BIn(wBMid16), .HiOut(wRegInB16), .LoOut(wRegInA17) );
BubbleSort_Node #( 32 ) BSN2_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid17), .BIn(wBMid17), .HiOut(wRegInB17), .LoOut(wRegInA18) );
BubbleSort_Node #( 32 ) BSN2_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid18), .BIn(wBMid18), .HiOut(wRegInB18), .LoOut(wRegInA19) );
BubbleSort_Node #( 32 ) BSN2_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid19), .BIn(wBMid19), .HiOut(wRegInB19), .LoOut(wRegInA20) );
BubbleSort_Node #( 32 ) BSN2_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid20), .BIn(wBMid20), .HiOut(wRegInB20), .LoOut(wRegInA21) );
BubbleSort_Node #( 32 ) BSN2_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid21), .BIn(wBMid21), .HiOut(wRegInB21), .LoOut(wRegInA22) );
BubbleSort_Node #( 32 ) BSN2_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid22), .BIn(wBMid22), .HiOut(wRegInB22), .LoOut(wRegInA23) );
BubbleSort_Node #( 32 ) BSN2_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid23), .BIn(wBMid23), .HiOut(wRegInB23), .LoOut(wRegInA24) );
BubbleSort_Node #( 32 ) BSN2_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid24), .BIn(wBMid24), .HiOut(wRegInB24), .LoOut(wRegInA25) );
BubbleSort_Node #( 32 ) BSN2_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid25), .BIn(wBMid25), .HiOut(wRegInB25), .LoOut(wRegInA26) );
BubbleSort_Node #( 32 ) BSN2_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid26), .BIn(wBMid26), .HiOut(wRegInB26), .LoOut(wRegInA27) );
BubbleSort_Node #( 32 ) BSN2_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid27), .BIn(wBMid27), .HiOut(wRegInB27), .LoOut(wRegInA28) );
BubbleSort_Node #( 32 ) BSN2_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid28), .BIn(wBMid28), .HiOut(wRegInB28), .LoOut(wRegInA29) );
BubbleSort_Node #( 32 ) BSN2_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid29), .BIn(wBMid29), .HiOut(wRegInB29), .LoOut(wRegInA30) );
BubbleSort_Node #( 32 ) BSN2_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid30), .BIn(wBMid30), .HiOut(wRegInB30), .LoOut(wRegInA31) );
BubbleSort_Node #( 32 ) BSN2_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid31), .BIn(wBMid31), .HiOut(wRegInB31), .LoOut(wRegInA32) );
BubbleSort_Node #( 32 ) BSN2_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid32), .BIn(wBMid32), .HiOut(wRegInB32), .LoOut(wRegInA33) );
BubbleSort_Node #( 32 ) BSN2_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid33), .BIn(wBMid33), .HiOut(wRegInB33), .LoOut(wRegInA34) );
BubbleSort_Node #( 32 ) BSN2_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid34), .BIn(wBMid34), .HiOut(wRegInB34), .LoOut(wRegInA35) );
BubbleSort_Node #( 32 ) BSN2_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid35), .BIn(wBMid35), .HiOut(wRegInB35), .LoOut(wRegInA36) );
BubbleSort_Node #( 32 ) BSN2_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid36), .BIn(wBMid36), .HiOut(wRegInB36), .LoOut(wRegInA37) );
BubbleSort_Node #( 32 ) BSN2_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid37), .BIn(wBMid37), .HiOut(wRegInB37), .LoOut(wRegInA38) );
BubbleSort_Node #( 32 ) BSN2_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid38), .BIn(wBMid38), .HiOut(wRegInB38), .LoOut(wRegInA39) );
BubbleSort_Node #( 32 ) BSN2_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid39), .BIn(wBMid39), .HiOut(wRegInB39), .LoOut(wRegInA40) );
BubbleSort_Node #( 32 ) BSN2_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid40), .BIn(wBMid40), .HiOut(wRegInB40), .LoOut(wRegInA41) );
BubbleSort_Node #( 32 ) BSN2_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid41), .BIn(wBMid41), .HiOut(wRegInB41), .LoOut(wRegInA42) );
BubbleSort_Node #( 32 ) BSN2_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid42), .BIn(wBMid42), .HiOut(wRegInB42), .LoOut(wRegInA43) );
BubbleSort_Node #( 32 ) BSN2_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid43), .BIn(wBMid43), .HiOut(wRegInB43), .LoOut(wRegInA44) );
BubbleSort_Node #( 32 ) BSN2_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid44), .BIn(wBMid44), .HiOut(wRegInB44), .LoOut(wRegInA45) );
BubbleSort_Node #( 32 ) BSN2_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid45), .BIn(wBMid45), .HiOut(wRegInB45), .LoOut(wRegInA46) );
BubbleSort_Node #( 32 ) BSN2_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid46), .BIn(wBMid46), .HiOut(wRegInB46), .LoOut(wRegInA47) );
BubbleSort_Node #( 32 ) BSN2_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid47), .BIn(wBMid47), .HiOut(wRegInB47), .LoOut(wRegInA48) );
BubbleSort_Node #( 32 ) BSN2_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid48), .BIn(wBMid48), .HiOut(wRegInB48), .LoOut(wRegInA49) );
BubbleSort_Node #( 32 ) BSN2_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid49), .BIn(wBMid49), .HiOut(wRegInB49), .LoOut(wRegInA50) );
BubbleSort_Node #( 32 ) BSN2_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid50), .BIn(wBMid50), .HiOut(wRegInB50), .LoOut(wRegInA51) );
BubbleSort_Node #( 32 ) BSN2_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid51), .BIn(wBMid51), .HiOut(wRegInB51), .LoOut(wRegInA52) );
BubbleSort_Node #( 32 ) BSN2_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid52), .BIn(wBMid52), .HiOut(wRegInB52), .LoOut(wRegInA53) );
BubbleSort_Node #( 32 ) BSN2_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid53), .BIn(wBMid53), .HiOut(wRegInB53), .LoOut(wRegInA54) );
BubbleSort_Node #( 32 ) BSN2_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid54), .BIn(wBMid54), .HiOut(wRegInB54), .LoOut(wRegInA55) );
BubbleSort_Node #( 32 ) BSN2_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid55), .BIn(wBMid55), .HiOut(wRegInB55), .LoOut(wRegInA56) );
BubbleSort_Node #( 32 ) BSN2_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid56), .BIn(wBMid56), .HiOut(wRegInB56), .LoOut(wRegInA57) );
BubbleSort_Node #( 32 ) BSN2_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid57), .BIn(wBMid57), .HiOut(wRegInB57), .LoOut(wRegInA58) );
BubbleSort_Node #( 32 ) BSN2_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid58), .BIn(wBMid58), .HiOut(wRegInB58), .LoOut(wRegInA59) );
BubbleSort_Node #( 32 ) BSN2_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid59), .BIn(wBMid59), .HiOut(wRegInB59), .LoOut(wRegInA60) );
BubbleSort_Node #( 32 ) BSN2_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid60), .BIn(wBMid60), .HiOut(wRegInB60), .LoOut(wRegInA61) );
BubbleSort_Node #( 32 ) BSN2_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid61), .BIn(wBMid61), .HiOut(wRegInB61), .LoOut(wRegInA62) );
BubbleSort_Node #( 32 ) BSN2_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid62), .BIn(wBMid62), .HiOut(wRegInB62), .LoOut(wRegInA63) );
BubbleSort_Node #( 32 ) BSN2_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid63), .BIn(wBMid63), .HiOut(wRegInB63), .LoOut(wRegInA64) );
BubbleSort_Node #( 32 ) BSN2_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid64), .BIn(wBMid64), .HiOut(wRegInB64), .LoOut(wRegInA65) );
BubbleSort_Node #( 32 ) BSN2_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid65), .BIn(wBMid65), .HiOut(wRegInB65), .LoOut(wRegInA66) );
BubbleSort_Node #( 32 ) BSN2_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid66), .BIn(wBMid66), .HiOut(wRegInB66), .LoOut(wRegInA67) );
BubbleSort_Node #( 32 ) BSN2_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid67), .BIn(wBMid67), .HiOut(wRegInB67), .LoOut(wRegInA68) );
BubbleSort_Node #( 32 ) BSN2_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid68), .BIn(wBMid68), .HiOut(wRegInB68), .LoOut(wRegInA69) );
BubbleSort_Node #( 32 ) BSN2_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid69), .BIn(wBMid69), .HiOut(wRegInB69), .LoOut(wRegInA70) );
BubbleSort_Node #( 32 ) BSN2_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid70), .BIn(wBMid70), .HiOut(wRegInB70), .LoOut(wRegInA71) );
BubbleSort_Node #( 32 ) BSN2_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid71), .BIn(wBMid71), .HiOut(wRegInB71), .LoOut(wRegInA72) );
BubbleSort_Node #( 32 ) BSN2_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid72), .BIn(wBMid72), .HiOut(wRegInB72), .LoOut(wRegInA73) );
BubbleSort_Node #( 32 ) BSN2_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid73), .BIn(wBMid73), .HiOut(wRegInB73), .LoOut(wRegInA74) );
BubbleSort_Node #( 32 ) BSN2_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid74), .BIn(wBMid74), .HiOut(wRegInB74), .LoOut(wRegInA75) );
BubbleSort_Node #( 32 ) BSN2_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid75), .BIn(wBMid75), .HiOut(wRegInB75), .LoOut(wRegInA76) );
BubbleSort_Node #( 32 ) BSN2_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid76), .BIn(wBMid76), .HiOut(wRegInB76), .LoOut(wRegInA77) );
BubbleSort_Node #( 32 ) BSN2_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid77), .BIn(wBMid77), .HiOut(wRegInB77), .LoOut(wRegInA78) );
BubbleSort_Node #( 32 ) BSN2_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid78), .BIn(wBMid78), .HiOut(wRegInB78), .LoOut(wRegInA79) );
BubbleSort_Node #( 32 ) BSN2_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid79), .BIn(wBMid79), .HiOut(wRegInB79), .LoOut(wRegInA80) );
BubbleSort_Node #( 32 ) BSN2_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid80), .BIn(wBMid80), .HiOut(wRegInB80), .LoOut(wRegInA81) );
BubbleSort_Node #( 32 ) BSN2_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid81), .BIn(wBMid81), .HiOut(wRegInB81), .LoOut(wRegInA82) );
BubbleSort_Node #( 32 ) BSN2_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid82), .BIn(wBMid82), .HiOut(wRegInB82), .LoOut(wRegInA83) );
BubbleSort_Node #( 32 ) BSN2_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid83), .BIn(wBMid83), .HiOut(wRegInB83), .LoOut(wRegInA84) );
BubbleSort_Node #( 32 ) BSN2_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid84), .BIn(wBMid84), .HiOut(wRegInB84), .LoOut(wRegInA85) );
BubbleSort_Node #( 32 ) BSN2_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid85), .BIn(wBMid85), .HiOut(wRegInB85), .LoOut(wRegInA86) );
BubbleSort_Node #( 32 ) BSN2_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid86), .BIn(wBMid86), .HiOut(wRegInB86), .LoOut(wRegInA87) );
BubbleSort_Node #( 32 ) BSN2_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid87), .BIn(wBMid87), .HiOut(wRegInB87), .LoOut(wRegInA88) );
BubbleSort_Node #( 32 ) BSN2_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid88), .BIn(wBMid88), .HiOut(wRegInB88), .LoOut(wRegInA89) );
BubbleSort_Node #( 32 ) BSN2_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid89), .BIn(wBMid89), .HiOut(wRegInB89), .LoOut(wRegInA90) );
BubbleSort_Node #( 32 ) BSN2_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid90), .BIn(wBMid90), .HiOut(wRegInB90), .LoOut(wRegInA91) );
BubbleSort_Node #( 32 ) BSN2_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid91), .BIn(wBMid91), .HiOut(wRegInB91), .LoOut(wRegInA92) );
BubbleSort_Node #( 32 ) BSN2_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid92), .BIn(wBMid92), .HiOut(wRegInB92), .LoOut(wRegInA93) );
BubbleSort_Node #( 32 ) BSN2_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid93), .BIn(wBMid93), .HiOut(wRegInB93), .LoOut(wRegInA94) );
BubbleSort_Node #( 32 ) BSN2_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid94), .BIn(wBMid94), .HiOut(wRegInB94), .LoOut(wRegInA95) );
BubbleSort_Node #( 32 ) BSN2_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid95), .BIn(wBMid95), .HiOut(wRegInB95), .LoOut(wRegInA96) );
BubbleSort_Node #( 32 ) BSN2_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid96), .BIn(wBMid96), .HiOut(wRegInB96), .LoOut(wRegInA97) );
BubbleSort_Node #( 32 ) BSN2_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid97), .BIn(wBMid97), .HiOut(wRegInB97), .LoOut(wRegInA98) );
BubbleSort_Node #( 32 ) BSN2_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid98), .BIn(wBMid98), .HiOut(wRegInB98), .LoOut(wRegInA99) );
BubbleSort_Node #( 32 ) BSN2_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid99), .BIn(wBMid99), .HiOut(wRegInB99), .LoOut(wRegInA100) );
BubbleSort_Node #( 32 ) BSN2_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid100), .BIn(wBMid100), .HiOut(wRegInB100), .LoOut(wRegInA101) );
BubbleSort_Node #( 32 ) BSN2_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid101), .BIn(wBMid101), .HiOut(wRegInB101), .LoOut(wRegInA102) );
BubbleSort_Node #( 32 ) BSN2_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid102), .BIn(wBMid102), .HiOut(wRegInB102), .LoOut(wRegInA103) );
BubbleSort_Node #( 32 ) BSN2_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid103), .BIn(wBMid103), .HiOut(wRegInB103), .LoOut(wRegInA104) );
BubbleSort_Node #( 32 ) BSN2_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid104), .BIn(wBMid104), .HiOut(wRegInB104), .LoOut(wRegInA105) );
BubbleSort_Node #( 32 ) BSN2_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid105), .BIn(wBMid105), .HiOut(wRegInB105), .LoOut(wRegInA106) );
BubbleSort_Node #( 32 ) BSN2_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid106), .BIn(wBMid106), .HiOut(wRegInB106), .LoOut(wRegInA107) );
BubbleSort_Node #( 32 ) BSN2_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid107), .BIn(wBMid107), .HiOut(wRegInB107), .LoOut(wRegInA108) );
BubbleSort_Node #( 32 ) BSN2_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid108), .BIn(wBMid108), .HiOut(wRegInB108), .LoOut(wRegInA109) );
BubbleSort_Node #( 32 ) BSN2_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid109), .BIn(wBMid109), .HiOut(wRegInB109), .LoOut(wRegInA110) );
BubbleSort_Node #( 32 ) BSN2_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid110), .BIn(wBMid110), .HiOut(wRegInB110), .LoOut(wRegInA111) );
BubbleSort_Node #( 32 ) BSN2_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid111), .BIn(wBMid111), .HiOut(wRegInB111), .LoOut(wRegInA112) );
BubbleSort_Node #( 32 ) BSN2_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid112), .BIn(wBMid112), .HiOut(wRegInB112), .LoOut(wRegInA113) );
BubbleSort_Node #( 32 ) BSN2_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid113), .BIn(wBMid113), .HiOut(wRegInB113), .LoOut(wRegInA114) );
BubbleSort_Node #( 32 ) BSN2_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid114), .BIn(wBMid114), .HiOut(wRegInB114), .LoOut(wRegInA115) );
BubbleSort_Node #( 32 ) BSN2_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid115), .BIn(wBMid115), .HiOut(wRegInB115), .LoOut(wRegInA116) );
BubbleSort_Node #( 32 ) BSN2_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid116), .BIn(wBMid116), .HiOut(wRegInB116), .LoOut(wRegInA117) );
BubbleSort_Node #( 32 ) BSN2_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid117), .BIn(wBMid117), .HiOut(wRegInB117), .LoOut(wRegInA118) );
BubbleSort_Node #( 32 ) BSN2_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid118), .BIn(wBMid118), .HiOut(wRegInB118), .LoOut(wRegInA119) );
BubbleSort_Node #( 32 ) BSN2_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid119), .BIn(wBMid119), .HiOut(wRegInB119), .LoOut(wRegInA120) );
BubbleSort_Node #( 32 ) BSN2_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid120), .BIn(wBMid120), .HiOut(wRegInB120), .LoOut(wRegInA121) );
BubbleSort_Node #( 32 ) BSN2_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid121), .BIn(wBMid121), .HiOut(wRegInB121), .LoOut(wRegInA122) );
BubbleSort_Node #( 32 ) BSN2_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid122), .BIn(wBMid122), .HiOut(wRegInB122), .LoOut(wRegInA123) );
BubbleSort_Node #( 32 ) BSN2_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid123), .BIn(wBMid123), .HiOut(wRegInB123), .LoOut(wRegInA124) );
BubbleSort_Node #( 32 ) BSN2_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid124), .BIn(wBMid124), .HiOut(wRegInB124), .LoOut(wRegInA125) );
BubbleSort_Node #( 32 ) BSN2_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid125), .BIn(wBMid125), .HiOut(wRegInB125), .LoOut(wRegInA126) );
BubbleSort_Node #( 32 ) BSN2_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid126), .BIn(wBMid126), .HiOut(wRegInB126), .LoOut(wRegInA127) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA0), .Out(wAIn0), .ScanIn(ScanLink256), .ScanOut(ScanLink255), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB0), .Out(wBIn0), .ScanIn(ScanLink255), .ScanOut(ScanLink254), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA1), .Out(wAIn1), .ScanIn(ScanLink254), .ScanOut(ScanLink253), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB1), .Out(wBIn1), .ScanIn(ScanLink253), .ScanOut(ScanLink252), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA2), .Out(wAIn2), .ScanIn(ScanLink252), .ScanOut(ScanLink251), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB2), .Out(wBIn2), .ScanIn(ScanLink251), .ScanOut(ScanLink250), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA3), .Out(wAIn3), .ScanIn(ScanLink250), .ScanOut(ScanLink249), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB3), .Out(wBIn3), .ScanIn(ScanLink249), .ScanOut(ScanLink248), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA4), .Out(wAIn4), .ScanIn(ScanLink248), .ScanOut(ScanLink247), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB4), .Out(wBIn4), .ScanIn(ScanLink247), .ScanOut(ScanLink246), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA5), .Out(wAIn5), .ScanIn(ScanLink246), .ScanOut(ScanLink245), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB5), .Out(wBIn5), .ScanIn(ScanLink245), .ScanOut(ScanLink244), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA6), .Out(wAIn6), .ScanIn(ScanLink244), .ScanOut(ScanLink243), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB6), .Out(wBIn6), .ScanIn(ScanLink243), .ScanOut(ScanLink242), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA7), .Out(wAIn7), .ScanIn(ScanLink242), .ScanOut(ScanLink241), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB7), .Out(wBIn7), .ScanIn(ScanLink241), .ScanOut(ScanLink240), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA8), .Out(wAIn8), .ScanIn(ScanLink240), .ScanOut(ScanLink239), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB8), .Out(wBIn8), .ScanIn(ScanLink239), .ScanOut(ScanLink238), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA9), .Out(wAIn9), .ScanIn(ScanLink238), .ScanOut(ScanLink237), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB9), .Out(wBIn9), .ScanIn(ScanLink237), .ScanOut(ScanLink236), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA10), .Out(wAIn10), .ScanIn(ScanLink236), .ScanOut(ScanLink235), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB10), .Out(wBIn10), .ScanIn(ScanLink235), .ScanOut(ScanLink234), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA11), .Out(wAIn11), .ScanIn(ScanLink234), .ScanOut(ScanLink233), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB11), .Out(wBIn11), .ScanIn(ScanLink233), .ScanOut(ScanLink232), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA12), .Out(wAIn12), .ScanIn(ScanLink232), .ScanOut(ScanLink231), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB12), .Out(wBIn12), .ScanIn(ScanLink231), .ScanOut(ScanLink230), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA13), .Out(wAIn13), .ScanIn(ScanLink230), .ScanOut(ScanLink229), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB13), .Out(wBIn13), .ScanIn(ScanLink229), .ScanOut(ScanLink228), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA14), .Out(wAIn14), .ScanIn(ScanLink228), .ScanOut(ScanLink227), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB14), .Out(wBIn14), .ScanIn(ScanLink227), .ScanOut(ScanLink226), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA15), .Out(wAIn15), .ScanIn(ScanLink226), .ScanOut(ScanLink225), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB15), .Out(wBIn15), .ScanIn(ScanLink225), .ScanOut(ScanLink224), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA16), .Out(wAIn16), .ScanIn(ScanLink224), .ScanOut(ScanLink223), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB16), .Out(wBIn16), .ScanIn(ScanLink223), .ScanOut(ScanLink222), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA17), .Out(wAIn17), .ScanIn(ScanLink222), .ScanOut(ScanLink221), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB17), .Out(wBIn17), .ScanIn(ScanLink221), .ScanOut(ScanLink220), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA18), .Out(wAIn18), .ScanIn(ScanLink220), .ScanOut(ScanLink219), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB18), .Out(wBIn18), .ScanIn(ScanLink219), .ScanOut(ScanLink218), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA19), .Out(wAIn19), .ScanIn(ScanLink218), .ScanOut(ScanLink217), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB19), .Out(wBIn19), .ScanIn(ScanLink217), .ScanOut(ScanLink216), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA20), .Out(wAIn20), .ScanIn(ScanLink216), .ScanOut(ScanLink215), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB20), .Out(wBIn20), .ScanIn(ScanLink215), .ScanOut(ScanLink214), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA21), .Out(wAIn21), .ScanIn(ScanLink214), .ScanOut(ScanLink213), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB21), .Out(wBIn21), .ScanIn(ScanLink213), .ScanOut(ScanLink212), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA22), .Out(wAIn22), .ScanIn(ScanLink212), .ScanOut(ScanLink211), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB22), .Out(wBIn22), .ScanIn(ScanLink211), .ScanOut(ScanLink210), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA23), .Out(wAIn23), .ScanIn(ScanLink210), .ScanOut(ScanLink209), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB23), .Out(wBIn23), .ScanIn(ScanLink209), .ScanOut(ScanLink208), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA24), .Out(wAIn24), .ScanIn(ScanLink208), .ScanOut(ScanLink207), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB24), .Out(wBIn24), .ScanIn(ScanLink207), .ScanOut(ScanLink206), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA25), .Out(wAIn25), .ScanIn(ScanLink206), .ScanOut(ScanLink205), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB25), .Out(wBIn25), .ScanIn(ScanLink205), .ScanOut(ScanLink204), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA26), .Out(wAIn26), .ScanIn(ScanLink204), .ScanOut(ScanLink203), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB26), .Out(wBIn26), .ScanIn(ScanLink203), .ScanOut(ScanLink202), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA27), .Out(wAIn27), .ScanIn(ScanLink202), .ScanOut(ScanLink201), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB27), .Out(wBIn27), .ScanIn(ScanLink201), .ScanOut(ScanLink200), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA28), .Out(wAIn28), .ScanIn(ScanLink200), .ScanOut(ScanLink199), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB28), .Out(wBIn28), .ScanIn(ScanLink199), .ScanOut(ScanLink198), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA29), .Out(wAIn29), .ScanIn(ScanLink198), .ScanOut(ScanLink197), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB29), .Out(wBIn29), .ScanIn(ScanLink197), .ScanOut(ScanLink196), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA30), .Out(wAIn30), .ScanIn(ScanLink196), .ScanOut(ScanLink195), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB30), .Out(wBIn30), .ScanIn(ScanLink195), .ScanOut(ScanLink194), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA31), .Out(wAIn31), .ScanIn(ScanLink194), .ScanOut(ScanLink193), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB31), .Out(wBIn31), .ScanIn(ScanLink193), .ScanOut(ScanLink192), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA32), .Out(wAIn32), .ScanIn(ScanLink192), .ScanOut(ScanLink191), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB32), .Out(wBIn32), .ScanIn(ScanLink191), .ScanOut(ScanLink190), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA33), .Out(wAIn33), .ScanIn(ScanLink190), .ScanOut(ScanLink189), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB33), .Out(wBIn33), .ScanIn(ScanLink189), .ScanOut(ScanLink188), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA34), .Out(wAIn34), .ScanIn(ScanLink188), .ScanOut(ScanLink187), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB34), .Out(wBIn34), .ScanIn(ScanLink187), .ScanOut(ScanLink186), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA35), .Out(wAIn35), .ScanIn(ScanLink186), .ScanOut(ScanLink185), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB35), .Out(wBIn35), .ScanIn(ScanLink185), .ScanOut(ScanLink184), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA36), .Out(wAIn36), .ScanIn(ScanLink184), .ScanOut(ScanLink183), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB36), .Out(wBIn36), .ScanIn(ScanLink183), .ScanOut(ScanLink182), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA37), .Out(wAIn37), .ScanIn(ScanLink182), .ScanOut(ScanLink181), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB37), .Out(wBIn37), .ScanIn(ScanLink181), .ScanOut(ScanLink180), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA38), .Out(wAIn38), .ScanIn(ScanLink180), .ScanOut(ScanLink179), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB38), .Out(wBIn38), .ScanIn(ScanLink179), .ScanOut(ScanLink178), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA39), .Out(wAIn39), .ScanIn(ScanLink178), .ScanOut(ScanLink177), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB39), .Out(wBIn39), .ScanIn(ScanLink177), .ScanOut(ScanLink176), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA40), .Out(wAIn40), .ScanIn(ScanLink176), .ScanOut(ScanLink175), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB40), .Out(wBIn40), .ScanIn(ScanLink175), .ScanOut(ScanLink174), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA41), .Out(wAIn41), .ScanIn(ScanLink174), .ScanOut(ScanLink173), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB41), .Out(wBIn41), .ScanIn(ScanLink173), .ScanOut(ScanLink172), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA42), .Out(wAIn42), .ScanIn(ScanLink172), .ScanOut(ScanLink171), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB42), .Out(wBIn42), .ScanIn(ScanLink171), .ScanOut(ScanLink170), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA43), .Out(wAIn43), .ScanIn(ScanLink170), .ScanOut(ScanLink169), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB43), .Out(wBIn43), .ScanIn(ScanLink169), .ScanOut(ScanLink168), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA44), .Out(wAIn44), .ScanIn(ScanLink168), .ScanOut(ScanLink167), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB44), .Out(wBIn44), .ScanIn(ScanLink167), .ScanOut(ScanLink166), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA45), .Out(wAIn45), .ScanIn(ScanLink166), .ScanOut(ScanLink165), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB45), .Out(wBIn45), .ScanIn(ScanLink165), .ScanOut(ScanLink164), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA46), .Out(wAIn46), .ScanIn(ScanLink164), .ScanOut(ScanLink163), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB46), .Out(wBIn46), .ScanIn(ScanLink163), .ScanOut(ScanLink162), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA47), .Out(wAIn47), .ScanIn(ScanLink162), .ScanOut(ScanLink161), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB47), .Out(wBIn47), .ScanIn(ScanLink161), .ScanOut(ScanLink160), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA48), .Out(wAIn48), .ScanIn(ScanLink160), .ScanOut(ScanLink159), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB48), .Out(wBIn48), .ScanIn(ScanLink159), .ScanOut(ScanLink158), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA49), .Out(wAIn49), .ScanIn(ScanLink158), .ScanOut(ScanLink157), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB49), .Out(wBIn49), .ScanIn(ScanLink157), .ScanOut(ScanLink156), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA50), .Out(wAIn50), .ScanIn(ScanLink156), .ScanOut(ScanLink155), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB50), .Out(wBIn50), .ScanIn(ScanLink155), .ScanOut(ScanLink154), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA51), .Out(wAIn51), .ScanIn(ScanLink154), .ScanOut(ScanLink153), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB51), .Out(wBIn51), .ScanIn(ScanLink153), .ScanOut(ScanLink152), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA52), .Out(wAIn52), .ScanIn(ScanLink152), .ScanOut(ScanLink151), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB52), .Out(wBIn52), .ScanIn(ScanLink151), .ScanOut(ScanLink150), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA53), .Out(wAIn53), .ScanIn(ScanLink150), .ScanOut(ScanLink149), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB53), .Out(wBIn53), .ScanIn(ScanLink149), .ScanOut(ScanLink148), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA54), .Out(wAIn54), .ScanIn(ScanLink148), .ScanOut(ScanLink147), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB54), .Out(wBIn54), .ScanIn(ScanLink147), .ScanOut(ScanLink146), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA55), .Out(wAIn55), .ScanIn(ScanLink146), .ScanOut(ScanLink145), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB55), .Out(wBIn55), .ScanIn(ScanLink145), .ScanOut(ScanLink144), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA56), .Out(wAIn56), .ScanIn(ScanLink144), .ScanOut(ScanLink143), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB56), .Out(wBIn56), .ScanIn(ScanLink143), .ScanOut(ScanLink142), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA57), .Out(wAIn57), .ScanIn(ScanLink142), .ScanOut(ScanLink141), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB57), .Out(wBIn57), .ScanIn(ScanLink141), .ScanOut(ScanLink140), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA58), .Out(wAIn58), .ScanIn(ScanLink140), .ScanOut(ScanLink139), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB58), .Out(wBIn58), .ScanIn(ScanLink139), .ScanOut(ScanLink138), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA59), .Out(wAIn59), .ScanIn(ScanLink138), .ScanOut(ScanLink137), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB59), .Out(wBIn59), .ScanIn(ScanLink137), .ScanOut(ScanLink136), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA60), .Out(wAIn60), .ScanIn(ScanLink136), .ScanOut(ScanLink135), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB60), .Out(wBIn60), .ScanIn(ScanLink135), .ScanOut(ScanLink134), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA61), .Out(wAIn61), .ScanIn(ScanLink134), .ScanOut(ScanLink133), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB61), .Out(wBIn61), .ScanIn(ScanLink133), .ScanOut(ScanLink132), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA62), .Out(wAIn62), .ScanIn(ScanLink132), .ScanOut(ScanLink131), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB62), .Out(wBIn62), .ScanIn(ScanLink131), .ScanOut(ScanLink130), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA63), .Out(wAIn63), .ScanIn(ScanLink130), .ScanOut(ScanLink129), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB63), .Out(wBIn63), .ScanIn(ScanLink129), .ScanOut(ScanLink128), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA64), .Out(wAIn64), .ScanIn(ScanLink128), .ScanOut(ScanLink127), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB64), .Out(wBIn64), .ScanIn(ScanLink127), .ScanOut(ScanLink126), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA65), .Out(wAIn65), .ScanIn(ScanLink126), .ScanOut(ScanLink125), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB65), .Out(wBIn65), .ScanIn(ScanLink125), .ScanOut(ScanLink124), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA66), .Out(wAIn66), .ScanIn(ScanLink124), .ScanOut(ScanLink123), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB66), .Out(wBIn66), .ScanIn(ScanLink123), .ScanOut(ScanLink122), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA67), .Out(wAIn67), .ScanIn(ScanLink122), .ScanOut(ScanLink121), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB67), .Out(wBIn67), .ScanIn(ScanLink121), .ScanOut(ScanLink120), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA68), .Out(wAIn68), .ScanIn(ScanLink120), .ScanOut(ScanLink119), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB68), .Out(wBIn68), .ScanIn(ScanLink119), .ScanOut(ScanLink118), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA69), .Out(wAIn69), .ScanIn(ScanLink118), .ScanOut(ScanLink117), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB69), .Out(wBIn69), .ScanIn(ScanLink117), .ScanOut(ScanLink116), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA70), .Out(wAIn70), .ScanIn(ScanLink116), .ScanOut(ScanLink115), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB70), .Out(wBIn70), .ScanIn(ScanLink115), .ScanOut(ScanLink114), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA71), .Out(wAIn71), .ScanIn(ScanLink114), .ScanOut(ScanLink113), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB71), .Out(wBIn71), .ScanIn(ScanLink113), .ScanOut(ScanLink112), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA72), .Out(wAIn72), .ScanIn(ScanLink112), .ScanOut(ScanLink111), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB72), .Out(wBIn72), .ScanIn(ScanLink111), .ScanOut(ScanLink110), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA73), .Out(wAIn73), .ScanIn(ScanLink110), .ScanOut(ScanLink109), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB73), .Out(wBIn73), .ScanIn(ScanLink109), .ScanOut(ScanLink108), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA74), .Out(wAIn74), .ScanIn(ScanLink108), .ScanOut(ScanLink107), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB74), .Out(wBIn74), .ScanIn(ScanLink107), .ScanOut(ScanLink106), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA75), .Out(wAIn75), .ScanIn(ScanLink106), .ScanOut(ScanLink105), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB75), .Out(wBIn75), .ScanIn(ScanLink105), .ScanOut(ScanLink104), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA76), .Out(wAIn76), .ScanIn(ScanLink104), .ScanOut(ScanLink103), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB76), .Out(wBIn76), .ScanIn(ScanLink103), .ScanOut(ScanLink102), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA77), .Out(wAIn77), .ScanIn(ScanLink102), .ScanOut(ScanLink101), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB77), .Out(wBIn77), .ScanIn(ScanLink101), .ScanOut(ScanLink100), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA78), .Out(wAIn78), .ScanIn(ScanLink100), .ScanOut(ScanLink99), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB78), .Out(wBIn78), .ScanIn(ScanLink99), .ScanOut(ScanLink98), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA79), .Out(wAIn79), .ScanIn(ScanLink98), .ScanOut(ScanLink97), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB79), .Out(wBIn79), .ScanIn(ScanLink97), .ScanOut(ScanLink96), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA80), .Out(wAIn80), .ScanIn(ScanLink96), .ScanOut(ScanLink95), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB80), .Out(wBIn80), .ScanIn(ScanLink95), .ScanOut(ScanLink94), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA81), .Out(wAIn81), .ScanIn(ScanLink94), .ScanOut(ScanLink93), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB81), .Out(wBIn81), .ScanIn(ScanLink93), .ScanOut(ScanLink92), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA82), .Out(wAIn82), .ScanIn(ScanLink92), .ScanOut(ScanLink91), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB82), .Out(wBIn82), .ScanIn(ScanLink91), .ScanOut(ScanLink90), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA83), .Out(wAIn83), .ScanIn(ScanLink90), .ScanOut(ScanLink89), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB83), .Out(wBIn83), .ScanIn(ScanLink89), .ScanOut(ScanLink88), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA84), .Out(wAIn84), .ScanIn(ScanLink88), .ScanOut(ScanLink87), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB84), .Out(wBIn84), .ScanIn(ScanLink87), .ScanOut(ScanLink86), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA85), .Out(wAIn85), .ScanIn(ScanLink86), .ScanOut(ScanLink85), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB85), .Out(wBIn85), .ScanIn(ScanLink85), .ScanOut(ScanLink84), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA86), .Out(wAIn86), .ScanIn(ScanLink84), .ScanOut(ScanLink83), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB86), .Out(wBIn86), .ScanIn(ScanLink83), .ScanOut(ScanLink82), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA87), .Out(wAIn87), .ScanIn(ScanLink82), .ScanOut(ScanLink81), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB87), .Out(wBIn87), .ScanIn(ScanLink81), .ScanOut(ScanLink80), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA88), .Out(wAIn88), .ScanIn(ScanLink80), .ScanOut(ScanLink79), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB88), .Out(wBIn88), .ScanIn(ScanLink79), .ScanOut(ScanLink78), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA89), .Out(wAIn89), .ScanIn(ScanLink78), .ScanOut(ScanLink77), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB89), .Out(wBIn89), .ScanIn(ScanLink77), .ScanOut(ScanLink76), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA90), .Out(wAIn90), .ScanIn(ScanLink76), .ScanOut(ScanLink75), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB90), .Out(wBIn90), .ScanIn(ScanLink75), .ScanOut(ScanLink74), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA91), .Out(wAIn91), .ScanIn(ScanLink74), .ScanOut(ScanLink73), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB91), .Out(wBIn91), .ScanIn(ScanLink73), .ScanOut(ScanLink72), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA92), .Out(wAIn92), .ScanIn(ScanLink72), .ScanOut(ScanLink71), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB92), .Out(wBIn92), .ScanIn(ScanLink71), .ScanOut(ScanLink70), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA93), .Out(wAIn93), .ScanIn(ScanLink70), .ScanOut(ScanLink69), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB93), .Out(wBIn93), .ScanIn(ScanLink69), .ScanOut(ScanLink68), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA94), .Out(wAIn94), .ScanIn(ScanLink68), .ScanOut(ScanLink67), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB94), .Out(wBIn94), .ScanIn(ScanLink67), .ScanOut(ScanLink66), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA95), .Out(wAIn95), .ScanIn(ScanLink66), .ScanOut(ScanLink65), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB95), .Out(wBIn95), .ScanIn(ScanLink65), .ScanOut(ScanLink64), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA96), .Out(wAIn96), .ScanIn(ScanLink64), .ScanOut(ScanLink63), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB96), .Out(wBIn96), .ScanIn(ScanLink63), .ScanOut(ScanLink62), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA97), .Out(wAIn97), .ScanIn(ScanLink62), .ScanOut(ScanLink61), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB97), .Out(wBIn97), .ScanIn(ScanLink61), .ScanOut(ScanLink60), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA98), .Out(wAIn98), .ScanIn(ScanLink60), .ScanOut(ScanLink59), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB98), .Out(wBIn98), .ScanIn(ScanLink59), .ScanOut(ScanLink58), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA99), .Out(wAIn99), .ScanIn(ScanLink58), .ScanOut(ScanLink57), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB99), .Out(wBIn99), .ScanIn(ScanLink57), .ScanOut(ScanLink56), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA100), .Out(wAIn100), .ScanIn(ScanLink56), .ScanOut(ScanLink55), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB100), .Out(wBIn100), .ScanIn(ScanLink55), .ScanOut(ScanLink54), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA101), .Out(wAIn101), .ScanIn(ScanLink54), .ScanOut(ScanLink53), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB101), .Out(wBIn101), .ScanIn(ScanLink53), .ScanOut(ScanLink52), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA102), .Out(wAIn102), .ScanIn(ScanLink52), .ScanOut(ScanLink51), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB102), .Out(wBIn102), .ScanIn(ScanLink51), .ScanOut(ScanLink50), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA103), .Out(wAIn103), .ScanIn(ScanLink50), .ScanOut(ScanLink49), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB103), .Out(wBIn103), .ScanIn(ScanLink49), .ScanOut(ScanLink48), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA104), .Out(wAIn104), .ScanIn(ScanLink48), .ScanOut(ScanLink47), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB104), .Out(wBIn104), .ScanIn(ScanLink47), .ScanOut(ScanLink46), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA105), .Out(wAIn105), .ScanIn(ScanLink46), .ScanOut(ScanLink45), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB105), .Out(wBIn105), .ScanIn(ScanLink45), .ScanOut(ScanLink44), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA106), .Out(wAIn106), .ScanIn(ScanLink44), .ScanOut(ScanLink43), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB106), .Out(wBIn106), .ScanIn(ScanLink43), .ScanOut(ScanLink42), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA107), .Out(wAIn107), .ScanIn(ScanLink42), .ScanOut(ScanLink41), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB107), .Out(wBIn107), .ScanIn(ScanLink41), .ScanOut(ScanLink40), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA108), .Out(wAIn108), .ScanIn(ScanLink40), .ScanOut(ScanLink39), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB108), .Out(wBIn108), .ScanIn(ScanLink39), .ScanOut(ScanLink38), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA109), .Out(wAIn109), .ScanIn(ScanLink38), .ScanOut(ScanLink37), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB109), .Out(wBIn109), .ScanIn(ScanLink37), .ScanOut(ScanLink36), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA110), .Out(wAIn110), .ScanIn(ScanLink36), .ScanOut(ScanLink35), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB110), .Out(wBIn110), .ScanIn(ScanLink35), .ScanOut(ScanLink34), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA111), .Out(wAIn111), .ScanIn(ScanLink34), .ScanOut(ScanLink33), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB111), .Out(wBIn111), .ScanIn(ScanLink33), .ScanOut(ScanLink32), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA112), .Out(wAIn112), .ScanIn(ScanLink32), .ScanOut(ScanLink31), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB112), .Out(wBIn112), .ScanIn(ScanLink31), .ScanOut(ScanLink30), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA113), .Out(wAIn113), .ScanIn(ScanLink30), .ScanOut(ScanLink29), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB113), .Out(wBIn113), .ScanIn(ScanLink29), .ScanOut(ScanLink28), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA114), .Out(wAIn114), .ScanIn(ScanLink28), .ScanOut(ScanLink27), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB114), .Out(wBIn114), .ScanIn(ScanLink27), .ScanOut(ScanLink26), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA115), .Out(wAIn115), .ScanIn(ScanLink26), .ScanOut(ScanLink25), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB115), .Out(wBIn115), .ScanIn(ScanLink25), .ScanOut(ScanLink24), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA116), .Out(wAIn116), .ScanIn(ScanLink24), .ScanOut(ScanLink23), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB116), .Out(wBIn116), .ScanIn(ScanLink23), .ScanOut(ScanLink22), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA117), .Out(wAIn117), .ScanIn(ScanLink22), .ScanOut(ScanLink21), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB117), .Out(wBIn117), .ScanIn(ScanLink21), .ScanOut(ScanLink20), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA118), .Out(wAIn118), .ScanIn(ScanLink20), .ScanOut(ScanLink19), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB118), .Out(wBIn118), .ScanIn(ScanLink19), .ScanOut(ScanLink18), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA119), .Out(wAIn119), .ScanIn(ScanLink18), .ScanOut(ScanLink17), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB119), .Out(wBIn119), .ScanIn(ScanLink17), .ScanOut(ScanLink16), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA120), .Out(wAIn120), .ScanIn(ScanLink16), .ScanOut(ScanLink15), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB120), .Out(wBIn120), .ScanIn(ScanLink15), .ScanOut(ScanLink14), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA121), .Out(wAIn121), .ScanIn(ScanLink14), .ScanOut(ScanLink13), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB121), .Out(wBIn121), .ScanIn(ScanLink13), .ScanOut(ScanLink12), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA122), .Out(wAIn122), .ScanIn(ScanLink12), .ScanOut(ScanLink11), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB122), .Out(wBIn122), .ScanIn(ScanLink11), .ScanOut(ScanLink10), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA123), .Out(wAIn123), .ScanIn(ScanLink10), .ScanOut(ScanLink9), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB123), .Out(wBIn123), .ScanIn(ScanLink9), .ScanOut(ScanLink8), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA124), .Out(wAIn124), .ScanIn(ScanLink8), .ScanOut(ScanLink7), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB124), .Out(wBIn124), .ScanIn(ScanLink7), .ScanOut(ScanLink6), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA125), .Out(wAIn125), .ScanIn(ScanLink6), .ScanOut(ScanLink5), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB125), .Out(wBIn125), .ScanIn(ScanLink5), .ScanOut(ScanLink4), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA126), .Out(wAIn126), .ScanIn(ScanLink4), .ScanOut(ScanLink3), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB126), .Out(wBIn126), .ScanIn(ScanLink3), .ScanOut(ScanLink2), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA127), .Out(wAIn127), .ScanIn(ScanLink2), .ScanOut(ScanLink1), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB127), .Out(wBIn127), .ScanIn(ScanLink1), .ScanOut(ScanLink0), .ScanEnable(ScanEnable) );
BubbleSort_Control #( 8, 1, 32, 1 ) U_BSC ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Enable(wEnable), .ScanIn(ScanLink0), .ScanOut(ScanLink256), .ScanEnable(ScanEnable), .ScanId(1'd0) );

/*
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
