

/*
 *
 * RAW Benchmark Suite main defines
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/bubblesort/src/library.v,v 1.4 1997/08/09 05:56:59 jbabb Exp $
 *
 * Library for Bubble Sort Benchmark
 *
 * Authors: Elliot Waingold         (elliotw@lcs.mit.edu)
 *          Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 BubbleSort_Node is the basic pairwise element comparator.  It
 outputs the greater of its two inputs to HiOut and the lower of
 the two to LoOut.
 */

module BubbleSort_Node (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
			AIn, BIn, HiOut, LoOut);

   parameter WIDTH = 8;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* local connections */

   input [WIDTH-1:0]		AIn, BIn;
   output [WIDTH-1:0]		HiOut, LoOut;
   wire				Predicate;

   assign Predicate = (AIn > BIn) ? 1 : 0;
   assign HiOut = (Predicate) ? AIn : BIn;
   assign LoOut = (Predicate) ? BIn : AIn;

endmodule


/*
 BubbleSort_Reg is a pipeline/input register that can be written
 to from the host interface as well as from its input wires.  It
 also has an enable input that must be high for it to clock data
 in from the inputs.
 */

module BubbleSort_Reg (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		       ScanIn, ScanOut, ScanEnable,
		       Id, Enable, In, Out);

   parameter			 WIDTH = 8,
				 IDWIDTH = 8,
				 SCAN = 1;

   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;


   /* local connections */

   input [IDWIDTH-1:0]		Id;
   input			Enable;
   input [WIDTH-1:0]		In;
   output [WIDTH-1:0]		Out;
   reg [WIDTH-1:0]		Out;


   /* support reading of the node data value (non-scan only) */

   assign DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out : `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;


   always @(posedge Clk)
      begin


	 /* reset will initialize the register to zero */

	 if (Reset)
	    Out = 0;


	 /* support scan in */

	 else if  (SCAN && ScanEnable)
	    Out = ScanIn[WIDTH-1:0];


	 /* support writing of the node data value (non-scan only) */

	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0] == Id))
	    Out = DataIn[WIDTH-1:0];

	 /* otherwise if enable is high, read in input data */

	 else if (Enable)
	    Out = In;

      end
endmodule


/*
 BubbleSort_Control is the control node.  When a value is written to
 it by the host, it holds the enable high for that number of clock
 periods.
 */

module BubbleSort_Control(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
			  ScanIn, ScanOut, ScanEnable, ScanId,
			  Id, Enable);

   parameter			 CWIDTH=8,
				 IDWIDTH=8,
				 WIDTH=8,
				 SCAN=1;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;
   input [IDWIDTH-1:0]		 ScanId;


   /* local connections */

   input [IDWIDTH-1:0]		 Id;
   output			 Enable;
   reg [CWIDTH-1:0]		 count;
   reg [WIDTH-1:0]		 ScanReg;


   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? count :
         (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;

   /* enable when count is active */

   assign Enable = !(count==0);


   always @(posedge Clk)
      begin


	 /* store current scan output */

	 ScanReg=ScanIn;


	 /* Logic to reset, write, and decrement the counter */

	 if (Reset)
	    count=0;
	 else if (WR && (Addr[IDWIDTH-1:0]==Id))
	    count=DataIn[CWIDTH-1:0];
	 else
	    if(count)
	       count=count-1;
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [31:0] wRegInA0;
wire [31:0] wRegInB0;
wire [31:0] wAIn0;
wire [31:0] wBIn0;
wire [31:0] wRegInA1;
wire [31:0] wRegInB1;
wire [31:0] wAIn1;
wire [31:0] wBIn1;
wire [31:0] wRegInA2;
wire [31:0] wRegInB2;
wire [31:0] wAIn2;
wire [31:0] wBIn2;
wire [31:0] wRegInA3;
wire [31:0] wRegInB3;
wire [31:0] wAIn3;
wire [31:0] wBIn3;
wire [31:0] wRegInA4;
wire [31:0] wRegInB4;
wire [31:0] wAIn4;
wire [31:0] wBIn4;
wire [31:0] wRegInA5;
wire [31:0] wRegInB5;
wire [31:0] wAIn5;
wire [31:0] wBIn5;
wire [31:0] wRegInA6;
wire [31:0] wRegInB6;
wire [31:0] wAIn6;
wire [31:0] wBIn6;
wire [31:0] wRegInA7;
wire [31:0] wRegInB7;
wire [31:0] wAIn7;
wire [31:0] wBIn7;
wire [31:0] wRegInA8;
wire [31:0] wRegInB8;
wire [31:0] wAIn8;
wire [31:0] wBIn8;
wire [31:0] wRegInA9;
wire [31:0] wRegInB9;
wire [31:0] wAIn9;
wire [31:0] wBIn9;
wire [31:0] wRegInA10;
wire [31:0] wRegInB10;
wire [31:0] wAIn10;
wire [31:0] wBIn10;
wire [31:0] wRegInA11;
wire [31:0] wRegInB11;
wire [31:0] wAIn11;
wire [31:0] wBIn11;
wire [31:0] wRegInA12;
wire [31:0] wRegInB12;
wire [31:0] wAIn12;
wire [31:0] wBIn12;
wire [31:0] wRegInA13;
wire [31:0] wRegInB13;
wire [31:0] wAIn13;
wire [31:0] wBIn13;
wire [31:0] wRegInA14;
wire [31:0] wRegInB14;
wire [31:0] wAIn14;
wire [31:0] wBIn14;
wire [31:0] wRegInA15;
wire [31:0] wRegInB15;
wire [31:0] wAIn15;
wire [31:0] wBIn15;
wire [31:0] wRegInA16;
wire [31:0] wRegInB16;
wire [31:0] wAIn16;
wire [31:0] wBIn16;
wire [31:0] wRegInA17;
wire [31:0] wRegInB17;
wire [31:0] wAIn17;
wire [31:0] wBIn17;
wire [31:0] wRegInA18;
wire [31:0] wRegInB18;
wire [31:0] wAIn18;
wire [31:0] wBIn18;
wire [31:0] wRegInA19;
wire [31:0] wRegInB19;
wire [31:0] wAIn19;
wire [31:0] wBIn19;
wire [31:0] wRegInA20;
wire [31:0] wRegInB20;
wire [31:0] wAIn20;
wire [31:0] wBIn20;
wire [31:0] wRegInA21;
wire [31:0] wRegInB21;
wire [31:0] wAIn21;
wire [31:0] wBIn21;
wire [31:0] wRegInA22;
wire [31:0] wRegInB22;
wire [31:0] wAIn22;
wire [31:0] wBIn22;
wire [31:0] wRegInA23;
wire [31:0] wRegInB23;
wire [31:0] wAIn23;
wire [31:0] wBIn23;
wire [31:0] wRegInA24;
wire [31:0] wRegInB24;
wire [31:0] wAIn24;
wire [31:0] wBIn24;
wire [31:0] wRegInA25;
wire [31:0] wRegInB25;
wire [31:0] wAIn25;
wire [31:0] wBIn25;
wire [31:0] wRegInA26;
wire [31:0] wRegInB26;
wire [31:0] wAIn26;
wire [31:0] wBIn26;
wire [31:0] wRegInA27;
wire [31:0] wRegInB27;
wire [31:0] wAIn27;
wire [31:0] wBIn27;
wire [31:0] wRegInA28;
wire [31:0] wRegInB28;
wire [31:0] wAIn28;
wire [31:0] wBIn28;
wire [31:0] wRegInA29;
wire [31:0] wRegInB29;
wire [31:0] wAIn29;
wire [31:0] wBIn29;
wire [31:0] wRegInA30;
wire [31:0] wRegInB30;
wire [31:0] wAIn30;
wire [31:0] wBIn30;
wire [31:0] wRegInA31;
wire [31:0] wRegInB31;
wire [31:0] wAIn31;
wire [31:0] wBIn31;
wire [31:0] wRegInA32;
wire [31:0] wRegInB32;
wire [31:0] wAIn32;
wire [31:0] wBIn32;
wire [31:0] wRegInA33;
wire [31:0] wRegInB33;
wire [31:0] wAIn33;
wire [31:0] wBIn33;
wire [31:0] wRegInA34;
wire [31:0] wRegInB34;
wire [31:0] wAIn34;
wire [31:0] wBIn34;
wire [31:0] wRegInA35;
wire [31:0] wRegInB35;
wire [31:0] wAIn35;
wire [31:0] wBIn35;
wire [31:0] wRegInA36;
wire [31:0] wRegInB36;
wire [31:0] wAIn36;
wire [31:0] wBIn36;
wire [31:0] wRegInA37;
wire [31:0] wRegInB37;
wire [31:0] wAIn37;
wire [31:0] wBIn37;
wire [31:0] wRegInA38;
wire [31:0] wRegInB38;
wire [31:0] wAIn38;
wire [31:0] wBIn38;
wire [31:0] wRegInA39;
wire [31:0] wRegInB39;
wire [31:0] wAIn39;
wire [31:0] wBIn39;
wire [31:0] wRegInA40;
wire [31:0] wRegInB40;
wire [31:0] wAIn40;
wire [31:0] wBIn40;
wire [31:0] wRegInA41;
wire [31:0] wRegInB41;
wire [31:0] wAIn41;
wire [31:0] wBIn41;
wire [31:0] wRegInA42;
wire [31:0] wRegInB42;
wire [31:0] wAIn42;
wire [31:0] wBIn42;
wire [31:0] wRegInA43;
wire [31:0] wRegInB43;
wire [31:0] wAIn43;
wire [31:0] wBIn43;
wire [31:0] wRegInA44;
wire [31:0] wRegInB44;
wire [31:0] wAIn44;
wire [31:0] wBIn44;
wire [31:0] wRegInA45;
wire [31:0] wRegInB45;
wire [31:0] wAIn45;
wire [31:0] wBIn45;
wire [31:0] wRegInA46;
wire [31:0] wRegInB46;
wire [31:0] wAIn46;
wire [31:0] wBIn46;
wire [31:0] wRegInA47;
wire [31:0] wRegInB47;
wire [31:0] wAIn47;
wire [31:0] wBIn47;
wire [31:0] wRegInA48;
wire [31:0] wRegInB48;
wire [31:0] wAIn48;
wire [31:0] wBIn48;
wire [31:0] wRegInA49;
wire [31:0] wRegInB49;
wire [31:0] wAIn49;
wire [31:0] wBIn49;
wire [31:0] wRegInA50;
wire [31:0] wRegInB50;
wire [31:0] wAIn50;
wire [31:0] wBIn50;
wire [31:0] wRegInA51;
wire [31:0] wRegInB51;
wire [31:0] wAIn51;
wire [31:0] wBIn51;
wire [31:0] wRegInA52;
wire [31:0] wRegInB52;
wire [31:0] wAIn52;
wire [31:0] wBIn52;
wire [31:0] wRegInA53;
wire [31:0] wRegInB53;
wire [31:0] wAIn53;
wire [31:0] wBIn53;
wire [31:0] wRegInA54;
wire [31:0] wRegInB54;
wire [31:0] wAIn54;
wire [31:0] wBIn54;
wire [31:0] wRegInA55;
wire [31:0] wRegInB55;
wire [31:0] wAIn55;
wire [31:0] wBIn55;
wire [31:0] wRegInA56;
wire [31:0] wRegInB56;
wire [31:0] wAIn56;
wire [31:0] wBIn56;
wire [31:0] wRegInA57;
wire [31:0] wRegInB57;
wire [31:0] wAIn57;
wire [31:0] wBIn57;
wire [31:0] wRegInA58;
wire [31:0] wRegInB58;
wire [31:0] wAIn58;
wire [31:0] wBIn58;
wire [31:0] wRegInA59;
wire [31:0] wRegInB59;
wire [31:0] wAIn59;
wire [31:0] wBIn59;
wire [31:0] wRegInA60;
wire [31:0] wRegInB60;
wire [31:0] wAIn60;
wire [31:0] wBIn60;
wire [31:0] wRegInA61;
wire [31:0] wRegInB61;
wire [31:0] wAIn61;
wire [31:0] wBIn61;
wire [31:0] wRegInA62;
wire [31:0] wRegInB62;
wire [31:0] wAIn62;
wire [31:0] wBIn62;
wire [31:0] wRegInA63;
wire [31:0] wRegInB63;
wire [31:0] wAIn63;
wire [31:0] wBIn63;
wire [31:0] wRegInA64;
wire [31:0] wRegInB64;
wire [31:0] wAIn64;
wire [31:0] wBIn64;
wire [31:0] wRegInA65;
wire [31:0] wRegInB65;
wire [31:0] wAIn65;
wire [31:0] wBIn65;
wire [31:0] wRegInA66;
wire [31:0] wRegInB66;
wire [31:0] wAIn66;
wire [31:0] wBIn66;
wire [31:0] wRegInA67;
wire [31:0] wRegInB67;
wire [31:0] wAIn67;
wire [31:0] wBIn67;
wire [31:0] wRegInA68;
wire [31:0] wRegInB68;
wire [31:0] wAIn68;
wire [31:0] wBIn68;
wire [31:0] wRegInA69;
wire [31:0] wRegInB69;
wire [31:0] wAIn69;
wire [31:0] wBIn69;
wire [31:0] wRegInA70;
wire [31:0] wRegInB70;
wire [31:0] wAIn70;
wire [31:0] wBIn70;
wire [31:0] wRegInA71;
wire [31:0] wRegInB71;
wire [31:0] wAIn71;
wire [31:0] wBIn71;
wire [31:0] wRegInA72;
wire [31:0] wRegInB72;
wire [31:0] wAIn72;
wire [31:0] wBIn72;
wire [31:0] wRegInA73;
wire [31:0] wRegInB73;
wire [31:0] wAIn73;
wire [31:0] wBIn73;
wire [31:0] wRegInA74;
wire [31:0] wRegInB74;
wire [31:0] wAIn74;
wire [31:0] wBIn74;
wire [31:0] wRegInA75;
wire [31:0] wRegInB75;
wire [31:0] wAIn75;
wire [31:0] wBIn75;
wire [31:0] wRegInA76;
wire [31:0] wRegInB76;
wire [31:0] wAIn76;
wire [31:0] wBIn76;
wire [31:0] wRegInA77;
wire [31:0] wRegInB77;
wire [31:0] wAIn77;
wire [31:0] wBIn77;
wire [31:0] wRegInA78;
wire [31:0] wRegInB78;
wire [31:0] wAIn78;
wire [31:0] wBIn78;
wire [31:0] wRegInA79;
wire [31:0] wRegInB79;
wire [31:0] wAIn79;
wire [31:0] wBIn79;
wire [31:0] wRegInA80;
wire [31:0] wRegInB80;
wire [31:0] wAIn80;
wire [31:0] wBIn80;
wire [31:0] wRegInA81;
wire [31:0] wRegInB81;
wire [31:0] wAIn81;
wire [31:0] wBIn81;
wire [31:0] wRegInA82;
wire [31:0] wRegInB82;
wire [31:0] wAIn82;
wire [31:0] wBIn82;
wire [31:0] wRegInA83;
wire [31:0] wRegInB83;
wire [31:0] wAIn83;
wire [31:0] wBIn83;
wire [31:0] wRegInA84;
wire [31:0] wRegInB84;
wire [31:0] wAIn84;
wire [31:0] wBIn84;
wire [31:0] wRegInA85;
wire [31:0] wRegInB85;
wire [31:0] wAIn85;
wire [31:0] wBIn85;
wire [31:0] wRegInA86;
wire [31:0] wRegInB86;
wire [31:0] wAIn86;
wire [31:0] wBIn86;
wire [31:0] wRegInA87;
wire [31:0] wRegInB87;
wire [31:0] wAIn87;
wire [31:0] wBIn87;
wire [31:0] wRegInA88;
wire [31:0] wRegInB88;
wire [31:0] wAIn88;
wire [31:0] wBIn88;
wire [31:0] wRegInA89;
wire [31:0] wRegInB89;
wire [31:0] wAIn89;
wire [31:0] wBIn89;
wire [31:0] wRegInA90;
wire [31:0] wRegInB90;
wire [31:0] wAIn90;
wire [31:0] wBIn90;
wire [31:0] wRegInA91;
wire [31:0] wRegInB91;
wire [31:0] wAIn91;
wire [31:0] wBIn91;
wire [31:0] wRegInA92;
wire [31:0] wRegInB92;
wire [31:0] wAIn92;
wire [31:0] wBIn92;
wire [31:0] wRegInA93;
wire [31:0] wRegInB93;
wire [31:0] wAIn93;
wire [31:0] wBIn93;
wire [31:0] wRegInA94;
wire [31:0] wRegInB94;
wire [31:0] wAIn94;
wire [31:0] wBIn94;
wire [31:0] wRegInA95;
wire [31:0] wRegInB95;
wire [31:0] wAIn95;
wire [31:0] wBIn95;
wire [31:0] wRegInA96;
wire [31:0] wRegInB96;
wire [31:0] wAIn96;
wire [31:0] wBIn96;
wire [31:0] wRegInA97;
wire [31:0] wRegInB97;
wire [31:0] wAIn97;
wire [31:0] wBIn97;
wire [31:0] wRegInA98;
wire [31:0] wRegInB98;
wire [31:0] wAIn98;
wire [31:0] wBIn98;
wire [31:0] wRegInA99;
wire [31:0] wRegInB99;
wire [31:0] wAIn99;
wire [31:0] wBIn99;
wire [31:0] wRegInA100;
wire [31:0] wRegInB100;
wire [31:0] wAIn100;
wire [31:0] wBIn100;
wire [31:0] wRegInA101;
wire [31:0] wRegInB101;
wire [31:0] wAIn101;
wire [31:0] wBIn101;
wire [31:0] wRegInA102;
wire [31:0] wRegInB102;
wire [31:0] wAIn102;
wire [31:0] wBIn102;
wire [31:0] wRegInA103;
wire [31:0] wRegInB103;
wire [31:0] wAIn103;
wire [31:0] wBIn103;
wire [31:0] wRegInA104;
wire [31:0] wRegInB104;
wire [31:0] wAIn104;
wire [31:0] wBIn104;
wire [31:0] wRegInA105;
wire [31:0] wRegInB105;
wire [31:0] wAIn105;
wire [31:0] wBIn105;
wire [31:0] wRegInA106;
wire [31:0] wRegInB106;
wire [31:0] wAIn106;
wire [31:0] wBIn106;
wire [31:0] wRegInA107;
wire [31:0] wRegInB107;
wire [31:0] wAIn107;
wire [31:0] wBIn107;
wire [31:0] wRegInA108;
wire [31:0] wRegInB108;
wire [31:0] wAIn108;
wire [31:0] wBIn108;
wire [31:0] wRegInA109;
wire [31:0] wRegInB109;
wire [31:0] wAIn109;
wire [31:0] wBIn109;
wire [31:0] wRegInA110;
wire [31:0] wRegInB110;
wire [31:0] wAIn110;
wire [31:0] wBIn110;
wire [31:0] wRegInA111;
wire [31:0] wRegInB111;
wire [31:0] wAIn111;
wire [31:0] wBIn111;
wire [31:0] wRegInA112;
wire [31:0] wRegInB112;
wire [31:0] wAIn112;
wire [31:0] wBIn112;
wire [31:0] wRegInA113;
wire [31:0] wRegInB113;
wire [31:0] wAIn113;
wire [31:0] wBIn113;
wire [31:0] wRegInA114;
wire [31:0] wRegInB114;
wire [31:0] wAIn114;
wire [31:0] wBIn114;
wire [31:0] wRegInA115;
wire [31:0] wRegInB115;
wire [31:0] wAIn115;
wire [31:0] wBIn115;
wire [31:0] wRegInA116;
wire [31:0] wRegInB116;
wire [31:0] wAIn116;
wire [31:0] wBIn116;
wire [31:0] wRegInA117;
wire [31:0] wRegInB117;
wire [31:0] wAIn117;
wire [31:0] wBIn117;
wire [31:0] wRegInA118;
wire [31:0] wRegInB118;
wire [31:0] wAIn118;
wire [31:0] wBIn118;
wire [31:0] wRegInA119;
wire [31:0] wRegInB119;
wire [31:0] wAIn119;
wire [31:0] wBIn119;
wire [31:0] wRegInA120;
wire [31:0] wRegInB120;
wire [31:0] wAIn120;
wire [31:0] wBIn120;
wire [31:0] wRegInA121;
wire [31:0] wRegInB121;
wire [31:0] wAIn121;
wire [31:0] wBIn121;
wire [31:0] wRegInA122;
wire [31:0] wRegInB122;
wire [31:0] wAIn122;
wire [31:0] wBIn122;
wire [31:0] wRegInA123;
wire [31:0] wRegInB123;
wire [31:0] wAIn123;
wire [31:0] wBIn123;
wire [31:0] wRegInA124;
wire [31:0] wRegInB124;
wire [31:0] wAIn124;
wire [31:0] wBIn124;
wire [31:0] wRegInA125;
wire [31:0] wRegInB125;
wire [31:0] wAIn125;
wire [31:0] wBIn125;
wire [31:0] wRegInA126;
wire [31:0] wRegInB126;
wire [31:0] wAIn126;
wire [31:0] wBIn126;
wire [31:0] wRegInA127;
wire [31:0] wRegInB127;
wire [31:0] wAIn127;
wire [31:0] wBIn127;
wire [31:0] wRegInA128;
wire [31:0] wRegInB128;
wire [31:0] wAIn128;
wire [31:0] wBIn128;
wire [31:0] wRegInA129;
wire [31:0] wRegInB129;
wire [31:0] wAIn129;
wire [31:0] wBIn129;
wire [31:0] wRegInA130;
wire [31:0] wRegInB130;
wire [31:0] wAIn130;
wire [31:0] wBIn130;
wire [31:0] wRegInA131;
wire [31:0] wRegInB131;
wire [31:0] wAIn131;
wire [31:0] wBIn131;
wire [31:0] wRegInA132;
wire [31:0] wRegInB132;
wire [31:0] wAIn132;
wire [31:0] wBIn132;
wire [31:0] wRegInA133;
wire [31:0] wRegInB133;
wire [31:0] wAIn133;
wire [31:0] wBIn133;
wire [31:0] wRegInA134;
wire [31:0] wRegInB134;
wire [31:0] wAIn134;
wire [31:0] wBIn134;
wire [31:0] wRegInA135;
wire [31:0] wRegInB135;
wire [31:0] wAIn135;
wire [31:0] wBIn135;
wire [31:0] wRegInA136;
wire [31:0] wRegInB136;
wire [31:0] wAIn136;
wire [31:0] wBIn136;
wire [31:0] wRegInA137;
wire [31:0] wRegInB137;
wire [31:0] wAIn137;
wire [31:0] wBIn137;
wire [31:0] wRegInA138;
wire [31:0] wRegInB138;
wire [31:0] wAIn138;
wire [31:0] wBIn138;
wire [31:0] wRegInA139;
wire [31:0] wRegInB139;
wire [31:0] wAIn139;
wire [31:0] wBIn139;
wire [31:0] wRegInA140;
wire [31:0] wRegInB140;
wire [31:0] wAIn140;
wire [31:0] wBIn140;
wire [31:0] wRegInA141;
wire [31:0] wRegInB141;
wire [31:0] wAIn141;
wire [31:0] wBIn141;
wire [31:0] wRegInA142;
wire [31:0] wRegInB142;
wire [31:0] wAIn142;
wire [31:0] wBIn142;
wire [31:0] wRegInA143;
wire [31:0] wRegInB143;
wire [31:0] wAIn143;
wire [31:0] wBIn143;
wire [31:0] wRegInA144;
wire [31:0] wRegInB144;
wire [31:0] wAIn144;
wire [31:0] wBIn144;
wire [31:0] wRegInA145;
wire [31:0] wRegInB145;
wire [31:0] wAIn145;
wire [31:0] wBIn145;
wire [31:0] wRegInA146;
wire [31:0] wRegInB146;
wire [31:0] wAIn146;
wire [31:0] wBIn146;
wire [31:0] wRegInA147;
wire [31:0] wRegInB147;
wire [31:0] wAIn147;
wire [31:0] wBIn147;
wire [31:0] wRegInA148;
wire [31:0] wRegInB148;
wire [31:0] wAIn148;
wire [31:0] wBIn148;
wire [31:0] wRegInA149;
wire [31:0] wRegInB149;
wire [31:0] wAIn149;
wire [31:0] wBIn149;
wire [31:0] wRegInA150;
wire [31:0] wRegInB150;
wire [31:0] wAIn150;
wire [31:0] wBIn150;
wire [31:0] wRegInA151;
wire [31:0] wRegInB151;
wire [31:0] wAIn151;
wire [31:0] wBIn151;
wire [31:0] wRegInA152;
wire [31:0] wRegInB152;
wire [31:0] wAIn152;
wire [31:0] wBIn152;
wire [31:0] wRegInA153;
wire [31:0] wRegInB153;
wire [31:0] wAIn153;
wire [31:0] wBIn153;
wire [31:0] wRegInA154;
wire [31:0] wRegInB154;
wire [31:0] wAIn154;
wire [31:0] wBIn154;
wire [31:0] wRegInA155;
wire [31:0] wRegInB155;
wire [31:0] wAIn155;
wire [31:0] wBIn155;
wire [31:0] wRegInA156;
wire [31:0] wRegInB156;
wire [31:0] wAIn156;
wire [31:0] wBIn156;
wire [31:0] wRegInA157;
wire [31:0] wRegInB157;
wire [31:0] wAIn157;
wire [31:0] wBIn157;
wire [31:0] wRegInA158;
wire [31:0] wRegInB158;
wire [31:0] wAIn158;
wire [31:0] wBIn158;
wire [31:0] wRegInA159;
wire [31:0] wRegInB159;
wire [31:0] wAIn159;
wire [31:0] wBIn159;
wire [31:0] wRegInA160;
wire [31:0] wRegInB160;
wire [31:0] wAIn160;
wire [31:0] wBIn160;
wire [31:0] wRegInA161;
wire [31:0] wRegInB161;
wire [31:0] wAIn161;
wire [31:0] wBIn161;
wire [31:0] wRegInA162;
wire [31:0] wRegInB162;
wire [31:0] wAIn162;
wire [31:0] wBIn162;
wire [31:0] wRegInA163;
wire [31:0] wRegInB163;
wire [31:0] wAIn163;
wire [31:0] wBIn163;
wire [31:0] wRegInA164;
wire [31:0] wRegInB164;
wire [31:0] wAIn164;
wire [31:0] wBIn164;
wire [31:0] wRegInA165;
wire [31:0] wRegInB165;
wire [31:0] wAIn165;
wire [31:0] wBIn165;
wire [31:0] wRegInA166;
wire [31:0] wRegInB166;
wire [31:0] wAIn166;
wire [31:0] wBIn166;
wire [31:0] wRegInA167;
wire [31:0] wRegInB167;
wire [31:0] wAIn167;
wire [31:0] wBIn167;
wire [31:0] wRegInA168;
wire [31:0] wRegInB168;
wire [31:0] wAIn168;
wire [31:0] wBIn168;
wire [31:0] wRegInA169;
wire [31:0] wRegInB169;
wire [31:0] wAIn169;
wire [31:0] wBIn169;
wire [31:0] wRegInA170;
wire [31:0] wRegInB170;
wire [31:0] wAIn170;
wire [31:0] wBIn170;
wire [31:0] wRegInA171;
wire [31:0] wRegInB171;
wire [31:0] wAIn171;
wire [31:0] wBIn171;
wire [31:0] wRegInA172;
wire [31:0] wRegInB172;
wire [31:0] wAIn172;
wire [31:0] wBIn172;
wire [31:0] wRegInA173;
wire [31:0] wRegInB173;
wire [31:0] wAIn173;
wire [31:0] wBIn173;
wire [31:0] wRegInA174;
wire [31:0] wRegInB174;
wire [31:0] wAIn174;
wire [31:0] wBIn174;
wire [31:0] wRegInA175;
wire [31:0] wRegInB175;
wire [31:0] wAIn175;
wire [31:0] wBIn175;
wire [31:0] wRegInA176;
wire [31:0] wRegInB176;
wire [31:0] wAIn176;
wire [31:0] wBIn176;
wire [31:0] wRegInA177;
wire [31:0] wRegInB177;
wire [31:0] wAIn177;
wire [31:0] wBIn177;
wire [31:0] wRegInA178;
wire [31:0] wRegInB178;
wire [31:0] wAIn178;
wire [31:0] wBIn178;
wire [31:0] wRegInA179;
wire [31:0] wRegInB179;
wire [31:0] wAIn179;
wire [31:0] wBIn179;
wire [31:0] wRegInA180;
wire [31:0] wRegInB180;
wire [31:0] wAIn180;
wire [31:0] wBIn180;
wire [31:0] wRegInA181;
wire [31:0] wRegInB181;
wire [31:0] wAIn181;
wire [31:0] wBIn181;
wire [31:0] wRegInA182;
wire [31:0] wRegInB182;
wire [31:0] wAIn182;
wire [31:0] wBIn182;
wire [31:0] wRegInA183;
wire [31:0] wRegInB183;
wire [31:0] wAIn183;
wire [31:0] wBIn183;
wire [31:0] wRegInA184;
wire [31:0] wRegInB184;
wire [31:0] wAIn184;
wire [31:0] wBIn184;
wire [31:0] wRegInA185;
wire [31:0] wRegInB185;
wire [31:0] wAIn185;
wire [31:0] wBIn185;
wire [31:0] wRegInA186;
wire [31:0] wRegInB186;
wire [31:0] wAIn186;
wire [31:0] wBIn186;
wire [31:0] wRegInA187;
wire [31:0] wRegInB187;
wire [31:0] wAIn187;
wire [31:0] wBIn187;
wire [31:0] wRegInA188;
wire [31:0] wRegInB188;
wire [31:0] wAIn188;
wire [31:0] wBIn188;
wire [31:0] wRegInA189;
wire [31:0] wRegInB189;
wire [31:0] wAIn189;
wire [31:0] wBIn189;
wire [31:0] wRegInA190;
wire [31:0] wRegInB190;
wire [31:0] wAIn190;
wire [31:0] wBIn190;
wire [31:0] wRegInA191;
wire [31:0] wRegInB191;
wire [31:0] wAIn191;
wire [31:0] wBIn191;
wire [31:0] wRegInA192;
wire [31:0] wRegInB192;
wire [31:0] wAIn192;
wire [31:0] wBIn192;
wire [31:0] wRegInA193;
wire [31:0] wRegInB193;
wire [31:0] wAIn193;
wire [31:0] wBIn193;
wire [31:0] wRegInA194;
wire [31:0] wRegInB194;
wire [31:0] wAIn194;
wire [31:0] wBIn194;
wire [31:0] wRegInA195;
wire [31:0] wRegInB195;
wire [31:0] wAIn195;
wire [31:0] wBIn195;
wire [31:0] wRegInA196;
wire [31:0] wRegInB196;
wire [31:0] wAIn196;
wire [31:0] wBIn196;
wire [31:0] wRegInA197;
wire [31:0] wRegInB197;
wire [31:0] wAIn197;
wire [31:0] wBIn197;
wire [31:0] wRegInA198;
wire [31:0] wRegInB198;
wire [31:0] wAIn198;
wire [31:0] wBIn198;
wire [31:0] wRegInA199;
wire [31:0] wRegInB199;
wire [31:0] wAIn199;
wire [31:0] wBIn199;
wire [31:0] wRegInA200;
wire [31:0] wRegInB200;
wire [31:0] wAIn200;
wire [31:0] wBIn200;
wire [31:0] wRegInA201;
wire [31:0] wRegInB201;
wire [31:0] wAIn201;
wire [31:0] wBIn201;
wire [31:0] wRegInA202;
wire [31:0] wRegInB202;
wire [31:0] wAIn202;
wire [31:0] wBIn202;
wire [31:0] wRegInA203;
wire [31:0] wRegInB203;
wire [31:0] wAIn203;
wire [31:0] wBIn203;
wire [31:0] wRegInA204;
wire [31:0] wRegInB204;
wire [31:0] wAIn204;
wire [31:0] wBIn204;
wire [31:0] wRegInA205;
wire [31:0] wRegInB205;
wire [31:0] wAIn205;
wire [31:0] wBIn205;
wire [31:0] wRegInA206;
wire [31:0] wRegInB206;
wire [31:0] wAIn206;
wire [31:0] wBIn206;
wire [31:0] wRegInA207;
wire [31:0] wRegInB207;
wire [31:0] wAIn207;
wire [31:0] wBIn207;
wire [31:0] wRegInA208;
wire [31:0] wRegInB208;
wire [31:0] wAIn208;
wire [31:0] wBIn208;
wire [31:0] wRegInA209;
wire [31:0] wRegInB209;
wire [31:0] wAIn209;
wire [31:0] wBIn209;
wire [31:0] wRegInA210;
wire [31:0] wRegInB210;
wire [31:0] wAIn210;
wire [31:0] wBIn210;
wire [31:0] wRegInA211;
wire [31:0] wRegInB211;
wire [31:0] wAIn211;
wire [31:0] wBIn211;
wire [31:0] wRegInA212;
wire [31:0] wRegInB212;
wire [31:0] wAIn212;
wire [31:0] wBIn212;
wire [31:0] wRegInA213;
wire [31:0] wRegInB213;
wire [31:0] wAIn213;
wire [31:0] wBIn213;
wire [31:0] wRegInA214;
wire [31:0] wRegInB214;
wire [31:0] wAIn214;
wire [31:0] wBIn214;
wire [31:0] wRegInA215;
wire [31:0] wRegInB215;
wire [31:0] wAIn215;
wire [31:0] wBIn215;
wire [31:0] wRegInA216;
wire [31:0] wRegInB216;
wire [31:0] wAIn216;
wire [31:0] wBIn216;
wire [31:0] wRegInA217;
wire [31:0] wRegInB217;
wire [31:0] wAIn217;
wire [31:0] wBIn217;
wire [31:0] wRegInA218;
wire [31:0] wRegInB218;
wire [31:0] wAIn218;
wire [31:0] wBIn218;
wire [31:0] wRegInA219;
wire [31:0] wRegInB219;
wire [31:0] wAIn219;
wire [31:0] wBIn219;
wire [31:0] wRegInA220;
wire [31:0] wRegInB220;
wire [31:0] wAIn220;
wire [31:0] wBIn220;
wire [31:0] wRegInA221;
wire [31:0] wRegInB221;
wire [31:0] wAIn221;
wire [31:0] wBIn221;
wire [31:0] wRegInA222;
wire [31:0] wRegInB222;
wire [31:0] wAIn222;
wire [31:0] wBIn222;
wire [31:0] wRegInA223;
wire [31:0] wRegInB223;
wire [31:0] wAIn223;
wire [31:0] wBIn223;
wire [31:0] wRegInA224;
wire [31:0] wRegInB224;
wire [31:0] wAIn224;
wire [31:0] wBIn224;
wire [31:0] wRegInA225;
wire [31:0] wRegInB225;
wire [31:0] wAIn225;
wire [31:0] wBIn225;
wire [31:0] wRegInA226;
wire [31:0] wRegInB226;
wire [31:0] wAIn226;
wire [31:0] wBIn226;
wire [31:0] wRegInA227;
wire [31:0] wRegInB227;
wire [31:0] wAIn227;
wire [31:0] wBIn227;
wire [31:0] wRegInA228;
wire [31:0] wRegInB228;
wire [31:0] wAIn228;
wire [31:0] wBIn228;
wire [31:0] wRegInA229;
wire [31:0] wRegInB229;
wire [31:0] wAIn229;
wire [31:0] wBIn229;
wire [31:0] wRegInA230;
wire [31:0] wRegInB230;
wire [31:0] wAIn230;
wire [31:0] wBIn230;
wire [31:0] wRegInA231;
wire [31:0] wRegInB231;
wire [31:0] wAIn231;
wire [31:0] wBIn231;
wire [31:0] wRegInA232;
wire [31:0] wRegInB232;
wire [31:0] wAIn232;
wire [31:0] wBIn232;
wire [31:0] wRegInA233;
wire [31:0] wRegInB233;
wire [31:0] wAIn233;
wire [31:0] wBIn233;
wire [31:0] wRegInA234;
wire [31:0] wRegInB234;
wire [31:0] wAIn234;
wire [31:0] wBIn234;
wire [31:0] wRegInA235;
wire [31:0] wRegInB235;
wire [31:0] wAIn235;
wire [31:0] wBIn235;
wire [31:0] wRegInA236;
wire [31:0] wRegInB236;
wire [31:0] wAIn236;
wire [31:0] wBIn236;
wire [31:0] wRegInA237;
wire [31:0] wRegInB237;
wire [31:0] wAIn237;
wire [31:0] wBIn237;
wire [31:0] wRegInA238;
wire [31:0] wRegInB238;
wire [31:0] wAIn238;
wire [31:0] wBIn238;
wire [31:0] wRegInA239;
wire [31:0] wRegInB239;
wire [31:0] wAIn239;
wire [31:0] wBIn239;
wire [31:0] wRegInA240;
wire [31:0] wRegInB240;
wire [31:0] wAIn240;
wire [31:0] wBIn240;
wire [31:0] wRegInA241;
wire [31:0] wRegInB241;
wire [31:0] wAIn241;
wire [31:0] wBIn241;
wire [31:0] wRegInA242;
wire [31:0] wRegInB242;
wire [31:0] wAIn242;
wire [31:0] wBIn242;
wire [31:0] wRegInA243;
wire [31:0] wRegInB243;
wire [31:0] wAIn243;
wire [31:0] wBIn243;
wire [31:0] wRegInA244;
wire [31:0] wRegInB244;
wire [31:0] wAIn244;
wire [31:0] wBIn244;
wire [31:0] wRegInA245;
wire [31:0] wRegInB245;
wire [31:0] wAIn245;
wire [31:0] wBIn245;
wire [31:0] wRegInA246;
wire [31:0] wRegInB246;
wire [31:0] wAIn246;
wire [31:0] wBIn246;
wire [31:0] wRegInA247;
wire [31:0] wRegInB247;
wire [31:0] wAIn247;
wire [31:0] wBIn247;
wire [31:0] wRegInA248;
wire [31:0] wRegInB248;
wire [31:0] wAIn248;
wire [31:0] wBIn248;
wire [31:0] wRegInA249;
wire [31:0] wRegInB249;
wire [31:0] wAIn249;
wire [31:0] wBIn249;
wire [31:0] wRegInA250;
wire [31:0] wRegInB250;
wire [31:0] wAIn250;
wire [31:0] wBIn250;
wire [31:0] wRegInA251;
wire [31:0] wRegInB251;
wire [31:0] wAIn251;
wire [31:0] wBIn251;
wire [31:0] wRegInA252;
wire [31:0] wRegInB252;
wire [31:0] wAIn252;
wire [31:0] wBIn252;
wire [31:0] wRegInA253;
wire [31:0] wRegInB253;
wire [31:0] wAIn253;
wire [31:0] wBIn253;
wire [31:0] wRegInA254;
wire [31:0] wRegInB254;
wire [31:0] wAIn254;
wire [31:0] wBIn254;
wire [31:0] wRegInA255;
wire [31:0] wRegInB255;
wire [31:0] wAIn255;
wire [31:0] wBIn255;
wire [31:0] wAMid0;
wire [31:0] wBMid0;
wire [31:0] wAMid1;
wire [31:0] wBMid1;
wire [31:0] wAMid2;
wire [31:0] wBMid2;
wire [31:0] wAMid3;
wire [31:0] wBMid3;
wire [31:0] wAMid4;
wire [31:0] wBMid4;
wire [31:0] wAMid5;
wire [31:0] wBMid5;
wire [31:0] wAMid6;
wire [31:0] wBMid6;
wire [31:0] wAMid7;
wire [31:0] wBMid7;
wire [31:0] wAMid8;
wire [31:0] wBMid8;
wire [31:0] wAMid9;
wire [31:0] wBMid9;
wire [31:0] wAMid10;
wire [31:0] wBMid10;
wire [31:0] wAMid11;
wire [31:0] wBMid11;
wire [31:0] wAMid12;
wire [31:0] wBMid12;
wire [31:0] wAMid13;
wire [31:0] wBMid13;
wire [31:0] wAMid14;
wire [31:0] wBMid14;
wire [31:0] wAMid15;
wire [31:0] wBMid15;
wire [31:0] wAMid16;
wire [31:0] wBMid16;
wire [31:0] wAMid17;
wire [31:0] wBMid17;
wire [31:0] wAMid18;
wire [31:0] wBMid18;
wire [31:0] wAMid19;
wire [31:0] wBMid19;
wire [31:0] wAMid20;
wire [31:0] wBMid20;
wire [31:0] wAMid21;
wire [31:0] wBMid21;
wire [31:0] wAMid22;
wire [31:0] wBMid22;
wire [31:0] wAMid23;
wire [31:0] wBMid23;
wire [31:0] wAMid24;
wire [31:0] wBMid24;
wire [31:0] wAMid25;
wire [31:0] wBMid25;
wire [31:0] wAMid26;
wire [31:0] wBMid26;
wire [31:0] wAMid27;
wire [31:0] wBMid27;
wire [31:0] wAMid28;
wire [31:0] wBMid28;
wire [31:0] wAMid29;
wire [31:0] wBMid29;
wire [31:0] wAMid30;
wire [31:0] wBMid30;
wire [31:0] wAMid31;
wire [31:0] wBMid31;
wire [31:0] wAMid32;
wire [31:0] wBMid32;
wire [31:0] wAMid33;
wire [31:0] wBMid33;
wire [31:0] wAMid34;
wire [31:0] wBMid34;
wire [31:0] wAMid35;
wire [31:0] wBMid35;
wire [31:0] wAMid36;
wire [31:0] wBMid36;
wire [31:0] wAMid37;
wire [31:0] wBMid37;
wire [31:0] wAMid38;
wire [31:0] wBMid38;
wire [31:0] wAMid39;
wire [31:0] wBMid39;
wire [31:0] wAMid40;
wire [31:0] wBMid40;
wire [31:0] wAMid41;
wire [31:0] wBMid41;
wire [31:0] wAMid42;
wire [31:0] wBMid42;
wire [31:0] wAMid43;
wire [31:0] wBMid43;
wire [31:0] wAMid44;
wire [31:0] wBMid44;
wire [31:0] wAMid45;
wire [31:0] wBMid45;
wire [31:0] wAMid46;
wire [31:0] wBMid46;
wire [31:0] wAMid47;
wire [31:0] wBMid47;
wire [31:0] wAMid48;
wire [31:0] wBMid48;
wire [31:0] wAMid49;
wire [31:0] wBMid49;
wire [31:0] wAMid50;
wire [31:0] wBMid50;
wire [31:0] wAMid51;
wire [31:0] wBMid51;
wire [31:0] wAMid52;
wire [31:0] wBMid52;
wire [31:0] wAMid53;
wire [31:0] wBMid53;
wire [31:0] wAMid54;
wire [31:0] wBMid54;
wire [31:0] wAMid55;
wire [31:0] wBMid55;
wire [31:0] wAMid56;
wire [31:0] wBMid56;
wire [31:0] wAMid57;
wire [31:0] wBMid57;
wire [31:0] wAMid58;
wire [31:0] wBMid58;
wire [31:0] wAMid59;
wire [31:0] wBMid59;
wire [31:0] wAMid60;
wire [31:0] wBMid60;
wire [31:0] wAMid61;
wire [31:0] wBMid61;
wire [31:0] wAMid62;
wire [31:0] wBMid62;
wire [31:0] wAMid63;
wire [31:0] wBMid63;
wire [31:0] wAMid64;
wire [31:0] wBMid64;
wire [31:0] wAMid65;
wire [31:0] wBMid65;
wire [31:0] wAMid66;
wire [31:0] wBMid66;
wire [31:0] wAMid67;
wire [31:0] wBMid67;
wire [31:0] wAMid68;
wire [31:0] wBMid68;
wire [31:0] wAMid69;
wire [31:0] wBMid69;
wire [31:0] wAMid70;
wire [31:0] wBMid70;
wire [31:0] wAMid71;
wire [31:0] wBMid71;
wire [31:0] wAMid72;
wire [31:0] wBMid72;
wire [31:0] wAMid73;
wire [31:0] wBMid73;
wire [31:0] wAMid74;
wire [31:0] wBMid74;
wire [31:0] wAMid75;
wire [31:0] wBMid75;
wire [31:0] wAMid76;
wire [31:0] wBMid76;
wire [31:0] wAMid77;
wire [31:0] wBMid77;
wire [31:0] wAMid78;
wire [31:0] wBMid78;
wire [31:0] wAMid79;
wire [31:0] wBMid79;
wire [31:0] wAMid80;
wire [31:0] wBMid80;
wire [31:0] wAMid81;
wire [31:0] wBMid81;
wire [31:0] wAMid82;
wire [31:0] wBMid82;
wire [31:0] wAMid83;
wire [31:0] wBMid83;
wire [31:0] wAMid84;
wire [31:0] wBMid84;
wire [31:0] wAMid85;
wire [31:0] wBMid85;
wire [31:0] wAMid86;
wire [31:0] wBMid86;
wire [31:0] wAMid87;
wire [31:0] wBMid87;
wire [31:0] wAMid88;
wire [31:0] wBMid88;
wire [31:0] wAMid89;
wire [31:0] wBMid89;
wire [31:0] wAMid90;
wire [31:0] wBMid90;
wire [31:0] wAMid91;
wire [31:0] wBMid91;
wire [31:0] wAMid92;
wire [31:0] wBMid92;
wire [31:0] wAMid93;
wire [31:0] wBMid93;
wire [31:0] wAMid94;
wire [31:0] wBMid94;
wire [31:0] wAMid95;
wire [31:0] wBMid95;
wire [31:0] wAMid96;
wire [31:0] wBMid96;
wire [31:0] wAMid97;
wire [31:0] wBMid97;
wire [31:0] wAMid98;
wire [31:0] wBMid98;
wire [31:0] wAMid99;
wire [31:0] wBMid99;
wire [31:0] wAMid100;
wire [31:0] wBMid100;
wire [31:0] wAMid101;
wire [31:0] wBMid101;
wire [31:0] wAMid102;
wire [31:0] wBMid102;
wire [31:0] wAMid103;
wire [31:0] wBMid103;
wire [31:0] wAMid104;
wire [31:0] wBMid104;
wire [31:0] wAMid105;
wire [31:0] wBMid105;
wire [31:0] wAMid106;
wire [31:0] wBMid106;
wire [31:0] wAMid107;
wire [31:0] wBMid107;
wire [31:0] wAMid108;
wire [31:0] wBMid108;
wire [31:0] wAMid109;
wire [31:0] wBMid109;
wire [31:0] wAMid110;
wire [31:0] wBMid110;
wire [31:0] wAMid111;
wire [31:0] wBMid111;
wire [31:0] wAMid112;
wire [31:0] wBMid112;
wire [31:0] wAMid113;
wire [31:0] wBMid113;
wire [31:0] wAMid114;
wire [31:0] wBMid114;
wire [31:0] wAMid115;
wire [31:0] wBMid115;
wire [31:0] wAMid116;
wire [31:0] wBMid116;
wire [31:0] wAMid117;
wire [31:0] wBMid117;
wire [31:0] wAMid118;
wire [31:0] wBMid118;
wire [31:0] wAMid119;
wire [31:0] wBMid119;
wire [31:0] wAMid120;
wire [31:0] wBMid120;
wire [31:0] wAMid121;
wire [31:0] wBMid121;
wire [31:0] wAMid122;
wire [31:0] wBMid122;
wire [31:0] wAMid123;
wire [31:0] wBMid123;
wire [31:0] wAMid124;
wire [31:0] wBMid124;
wire [31:0] wAMid125;
wire [31:0] wBMid125;
wire [31:0] wAMid126;
wire [31:0] wBMid126;
wire [31:0] wAMid127;
wire [31:0] wBMid127;
wire [31:0] wAMid128;
wire [31:0] wBMid128;
wire [31:0] wAMid129;
wire [31:0] wBMid129;
wire [31:0] wAMid130;
wire [31:0] wBMid130;
wire [31:0] wAMid131;
wire [31:0] wBMid131;
wire [31:0] wAMid132;
wire [31:0] wBMid132;
wire [31:0] wAMid133;
wire [31:0] wBMid133;
wire [31:0] wAMid134;
wire [31:0] wBMid134;
wire [31:0] wAMid135;
wire [31:0] wBMid135;
wire [31:0] wAMid136;
wire [31:0] wBMid136;
wire [31:0] wAMid137;
wire [31:0] wBMid137;
wire [31:0] wAMid138;
wire [31:0] wBMid138;
wire [31:0] wAMid139;
wire [31:0] wBMid139;
wire [31:0] wAMid140;
wire [31:0] wBMid140;
wire [31:0] wAMid141;
wire [31:0] wBMid141;
wire [31:0] wAMid142;
wire [31:0] wBMid142;
wire [31:0] wAMid143;
wire [31:0] wBMid143;
wire [31:0] wAMid144;
wire [31:0] wBMid144;
wire [31:0] wAMid145;
wire [31:0] wBMid145;
wire [31:0] wAMid146;
wire [31:0] wBMid146;
wire [31:0] wAMid147;
wire [31:0] wBMid147;
wire [31:0] wAMid148;
wire [31:0] wBMid148;
wire [31:0] wAMid149;
wire [31:0] wBMid149;
wire [31:0] wAMid150;
wire [31:0] wBMid150;
wire [31:0] wAMid151;
wire [31:0] wBMid151;
wire [31:0] wAMid152;
wire [31:0] wBMid152;
wire [31:0] wAMid153;
wire [31:0] wBMid153;
wire [31:0] wAMid154;
wire [31:0] wBMid154;
wire [31:0] wAMid155;
wire [31:0] wBMid155;
wire [31:0] wAMid156;
wire [31:0] wBMid156;
wire [31:0] wAMid157;
wire [31:0] wBMid157;
wire [31:0] wAMid158;
wire [31:0] wBMid158;
wire [31:0] wAMid159;
wire [31:0] wBMid159;
wire [31:0] wAMid160;
wire [31:0] wBMid160;
wire [31:0] wAMid161;
wire [31:0] wBMid161;
wire [31:0] wAMid162;
wire [31:0] wBMid162;
wire [31:0] wAMid163;
wire [31:0] wBMid163;
wire [31:0] wAMid164;
wire [31:0] wBMid164;
wire [31:0] wAMid165;
wire [31:0] wBMid165;
wire [31:0] wAMid166;
wire [31:0] wBMid166;
wire [31:0] wAMid167;
wire [31:0] wBMid167;
wire [31:0] wAMid168;
wire [31:0] wBMid168;
wire [31:0] wAMid169;
wire [31:0] wBMid169;
wire [31:0] wAMid170;
wire [31:0] wBMid170;
wire [31:0] wAMid171;
wire [31:0] wBMid171;
wire [31:0] wAMid172;
wire [31:0] wBMid172;
wire [31:0] wAMid173;
wire [31:0] wBMid173;
wire [31:0] wAMid174;
wire [31:0] wBMid174;
wire [31:0] wAMid175;
wire [31:0] wBMid175;
wire [31:0] wAMid176;
wire [31:0] wBMid176;
wire [31:0] wAMid177;
wire [31:0] wBMid177;
wire [31:0] wAMid178;
wire [31:0] wBMid178;
wire [31:0] wAMid179;
wire [31:0] wBMid179;
wire [31:0] wAMid180;
wire [31:0] wBMid180;
wire [31:0] wAMid181;
wire [31:0] wBMid181;
wire [31:0] wAMid182;
wire [31:0] wBMid182;
wire [31:0] wAMid183;
wire [31:0] wBMid183;
wire [31:0] wAMid184;
wire [31:0] wBMid184;
wire [31:0] wAMid185;
wire [31:0] wBMid185;
wire [31:0] wAMid186;
wire [31:0] wBMid186;
wire [31:0] wAMid187;
wire [31:0] wBMid187;
wire [31:0] wAMid188;
wire [31:0] wBMid188;
wire [31:0] wAMid189;
wire [31:0] wBMid189;
wire [31:0] wAMid190;
wire [31:0] wBMid190;
wire [31:0] wAMid191;
wire [31:0] wBMid191;
wire [31:0] wAMid192;
wire [31:0] wBMid192;
wire [31:0] wAMid193;
wire [31:0] wBMid193;
wire [31:0] wAMid194;
wire [31:0] wBMid194;
wire [31:0] wAMid195;
wire [31:0] wBMid195;
wire [31:0] wAMid196;
wire [31:0] wBMid196;
wire [31:0] wAMid197;
wire [31:0] wBMid197;
wire [31:0] wAMid198;
wire [31:0] wBMid198;
wire [31:0] wAMid199;
wire [31:0] wBMid199;
wire [31:0] wAMid200;
wire [31:0] wBMid200;
wire [31:0] wAMid201;
wire [31:0] wBMid201;
wire [31:0] wAMid202;
wire [31:0] wBMid202;
wire [31:0] wAMid203;
wire [31:0] wBMid203;
wire [31:0] wAMid204;
wire [31:0] wBMid204;
wire [31:0] wAMid205;
wire [31:0] wBMid205;
wire [31:0] wAMid206;
wire [31:0] wBMid206;
wire [31:0] wAMid207;
wire [31:0] wBMid207;
wire [31:0] wAMid208;
wire [31:0] wBMid208;
wire [31:0] wAMid209;
wire [31:0] wBMid209;
wire [31:0] wAMid210;
wire [31:0] wBMid210;
wire [31:0] wAMid211;
wire [31:0] wBMid211;
wire [31:0] wAMid212;
wire [31:0] wBMid212;
wire [31:0] wAMid213;
wire [31:0] wBMid213;
wire [31:0] wAMid214;
wire [31:0] wBMid214;
wire [31:0] wAMid215;
wire [31:0] wBMid215;
wire [31:0] wAMid216;
wire [31:0] wBMid216;
wire [31:0] wAMid217;
wire [31:0] wBMid217;
wire [31:0] wAMid218;
wire [31:0] wBMid218;
wire [31:0] wAMid219;
wire [31:0] wBMid219;
wire [31:0] wAMid220;
wire [31:0] wBMid220;
wire [31:0] wAMid221;
wire [31:0] wBMid221;
wire [31:0] wAMid222;
wire [31:0] wBMid222;
wire [31:0] wAMid223;
wire [31:0] wBMid223;
wire [31:0] wAMid224;
wire [31:0] wBMid224;
wire [31:0] wAMid225;
wire [31:0] wBMid225;
wire [31:0] wAMid226;
wire [31:0] wBMid226;
wire [31:0] wAMid227;
wire [31:0] wBMid227;
wire [31:0] wAMid228;
wire [31:0] wBMid228;
wire [31:0] wAMid229;
wire [31:0] wBMid229;
wire [31:0] wAMid230;
wire [31:0] wBMid230;
wire [31:0] wAMid231;
wire [31:0] wBMid231;
wire [31:0] wAMid232;
wire [31:0] wBMid232;
wire [31:0] wAMid233;
wire [31:0] wBMid233;
wire [31:0] wAMid234;
wire [31:0] wBMid234;
wire [31:0] wAMid235;
wire [31:0] wBMid235;
wire [31:0] wAMid236;
wire [31:0] wBMid236;
wire [31:0] wAMid237;
wire [31:0] wBMid237;
wire [31:0] wAMid238;
wire [31:0] wBMid238;
wire [31:0] wAMid239;
wire [31:0] wBMid239;
wire [31:0] wAMid240;
wire [31:0] wBMid240;
wire [31:0] wAMid241;
wire [31:0] wBMid241;
wire [31:0] wAMid242;
wire [31:0] wBMid242;
wire [31:0] wAMid243;
wire [31:0] wBMid243;
wire [31:0] wAMid244;
wire [31:0] wBMid244;
wire [31:0] wAMid245;
wire [31:0] wBMid245;
wire [31:0] wAMid246;
wire [31:0] wBMid246;
wire [31:0] wAMid247;
wire [31:0] wBMid247;
wire [31:0] wAMid248;
wire [31:0] wBMid248;
wire [31:0] wAMid249;
wire [31:0] wBMid249;
wire [31:0] wAMid250;
wire [31:0] wBMid250;
wire [31:0] wAMid251;
wire [31:0] wBMid251;
wire [31:0] wAMid252;
wire [31:0] wBMid252;
wire [31:0] wAMid253;
wire [31:0] wBMid253;
wire [31:0] wAMid254;
wire [31:0] wBMid254;
wire [0:0] wEnable;
wire [0:0] ScanEnable;
wire [31:0] ScanLink0;
wire [31:0] ScanLink1;
wire [31:0] ScanLink2;
wire [31:0] ScanLink3;
wire [31:0] ScanLink4;
wire [31:0] ScanLink5;
wire [31:0] ScanLink6;
wire [31:0] ScanLink7;
wire [31:0] ScanLink8;
wire [31:0] ScanLink9;
wire [31:0] ScanLink10;
wire [31:0] ScanLink11;
wire [31:0] ScanLink12;
wire [31:0] ScanLink13;
wire [31:0] ScanLink14;
wire [31:0] ScanLink15;
wire [31:0] ScanLink16;
wire [31:0] ScanLink17;
wire [31:0] ScanLink18;
wire [31:0] ScanLink19;
wire [31:0] ScanLink20;
wire [31:0] ScanLink21;
wire [31:0] ScanLink22;
wire [31:0] ScanLink23;
wire [31:0] ScanLink24;
wire [31:0] ScanLink25;
wire [31:0] ScanLink26;
wire [31:0] ScanLink27;
wire [31:0] ScanLink28;
wire [31:0] ScanLink29;
wire [31:0] ScanLink30;
wire [31:0] ScanLink31;
wire [31:0] ScanLink32;
wire [31:0] ScanLink33;
wire [31:0] ScanLink34;
wire [31:0] ScanLink35;
wire [31:0] ScanLink36;
wire [31:0] ScanLink37;
wire [31:0] ScanLink38;
wire [31:0] ScanLink39;
wire [31:0] ScanLink40;
wire [31:0] ScanLink41;
wire [31:0] ScanLink42;
wire [31:0] ScanLink43;
wire [31:0] ScanLink44;
wire [31:0] ScanLink45;
wire [31:0] ScanLink46;
wire [31:0] ScanLink47;
wire [31:0] ScanLink48;
wire [31:0] ScanLink49;
wire [31:0] ScanLink50;
wire [31:0] ScanLink51;
wire [31:0] ScanLink52;
wire [31:0] ScanLink53;
wire [31:0] ScanLink54;
wire [31:0] ScanLink55;
wire [31:0] ScanLink56;
wire [31:0] ScanLink57;
wire [31:0] ScanLink58;
wire [31:0] ScanLink59;
wire [31:0] ScanLink60;
wire [31:0] ScanLink61;
wire [31:0] ScanLink62;
wire [31:0] ScanLink63;
wire [31:0] ScanLink64;
wire [31:0] ScanLink65;
wire [31:0] ScanLink66;
wire [31:0] ScanLink67;
wire [31:0] ScanLink68;
wire [31:0] ScanLink69;
wire [31:0] ScanLink70;
wire [31:0] ScanLink71;
wire [31:0] ScanLink72;
wire [31:0] ScanLink73;
wire [31:0] ScanLink74;
wire [31:0] ScanLink75;
wire [31:0] ScanLink76;
wire [31:0] ScanLink77;
wire [31:0] ScanLink78;
wire [31:0] ScanLink79;
wire [31:0] ScanLink80;
wire [31:0] ScanLink81;
wire [31:0] ScanLink82;
wire [31:0] ScanLink83;
wire [31:0] ScanLink84;
wire [31:0] ScanLink85;
wire [31:0] ScanLink86;
wire [31:0] ScanLink87;
wire [31:0] ScanLink88;
wire [31:0] ScanLink89;
wire [31:0] ScanLink90;
wire [31:0] ScanLink91;
wire [31:0] ScanLink92;
wire [31:0] ScanLink93;
wire [31:0] ScanLink94;
wire [31:0] ScanLink95;
wire [31:0] ScanLink96;
wire [31:0] ScanLink97;
wire [31:0] ScanLink98;
wire [31:0] ScanLink99;
wire [31:0] ScanLink100;
wire [31:0] ScanLink101;
wire [31:0] ScanLink102;
wire [31:0] ScanLink103;
wire [31:0] ScanLink104;
wire [31:0] ScanLink105;
wire [31:0] ScanLink106;
wire [31:0] ScanLink107;
wire [31:0] ScanLink108;
wire [31:0] ScanLink109;
wire [31:0] ScanLink110;
wire [31:0] ScanLink111;
wire [31:0] ScanLink112;
wire [31:0] ScanLink113;
wire [31:0] ScanLink114;
wire [31:0] ScanLink115;
wire [31:0] ScanLink116;
wire [31:0] ScanLink117;
wire [31:0] ScanLink118;
wire [31:0] ScanLink119;
wire [31:0] ScanLink120;
wire [31:0] ScanLink121;
wire [31:0] ScanLink122;
wire [31:0] ScanLink123;
wire [31:0] ScanLink124;
wire [31:0] ScanLink125;
wire [31:0] ScanLink126;
wire [31:0] ScanLink127;
wire [31:0] ScanLink128;
wire [31:0] ScanLink129;
wire [31:0] ScanLink130;
wire [31:0] ScanLink131;
wire [31:0] ScanLink132;
wire [31:0] ScanLink133;
wire [31:0] ScanLink134;
wire [31:0] ScanLink135;
wire [31:0] ScanLink136;
wire [31:0] ScanLink137;
wire [31:0] ScanLink138;
wire [31:0] ScanLink139;
wire [31:0] ScanLink140;
wire [31:0] ScanLink141;
wire [31:0] ScanLink142;
wire [31:0] ScanLink143;
wire [31:0] ScanLink144;
wire [31:0] ScanLink145;
wire [31:0] ScanLink146;
wire [31:0] ScanLink147;
wire [31:0] ScanLink148;
wire [31:0] ScanLink149;
wire [31:0] ScanLink150;
wire [31:0] ScanLink151;
wire [31:0] ScanLink152;
wire [31:0] ScanLink153;
wire [31:0] ScanLink154;
wire [31:0] ScanLink155;
wire [31:0] ScanLink156;
wire [31:0] ScanLink157;
wire [31:0] ScanLink158;
wire [31:0] ScanLink159;
wire [31:0] ScanLink160;
wire [31:0] ScanLink161;
wire [31:0] ScanLink162;
wire [31:0] ScanLink163;
wire [31:0] ScanLink164;
wire [31:0] ScanLink165;
wire [31:0] ScanLink166;
wire [31:0] ScanLink167;
wire [31:0] ScanLink168;
wire [31:0] ScanLink169;
wire [31:0] ScanLink170;
wire [31:0] ScanLink171;
wire [31:0] ScanLink172;
wire [31:0] ScanLink173;
wire [31:0] ScanLink174;
wire [31:0] ScanLink175;
wire [31:0] ScanLink176;
wire [31:0] ScanLink177;
wire [31:0] ScanLink178;
wire [31:0] ScanLink179;
wire [31:0] ScanLink180;
wire [31:0] ScanLink181;
wire [31:0] ScanLink182;
wire [31:0] ScanLink183;
wire [31:0] ScanLink184;
wire [31:0] ScanLink185;
wire [31:0] ScanLink186;
wire [31:0] ScanLink187;
wire [31:0] ScanLink188;
wire [31:0] ScanLink189;
wire [31:0] ScanLink190;
wire [31:0] ScanLink191;
wire [31:0] ScanLink192;
wire [31:0] ScanLink193;
wire [31:0] ScanLink194;
wire [31:0] ScanLink195;
wire [31:0] ScanLink196;
wire [31:0] ScanLink197;
wire [31:0] ScanLink198;
wire [31:0] ScanLink199;
wire [31:0] ScanLink200;
wire [31:0] ScanLink201;
wire [31:0] ScanLink202;
wire [31:0] ScanLink203;
wire [31:0] ScanLink204;
wire [31:0] ScanLink205;
wire [31:0] ScanLink206;
wire [31:0] ScanLink207;
wire [31:0] ScanLink208;
wire [31:0] ScanLink209;
wire [31:0] ScanLink210;
wire [31:0] ScanLink211;
wire [31:0] ScanLink212;
wire [31:0] ScanLink213;
wire [31:0] ScanLink214;
wire [31:0] ScanLink215;
wire [31:0] ScanLink216;
wire [31:0] ScanLink217;
wire [31:0] ScanLink218;
wire [31:0] ScanLink219;
wire [31:0] ScanLink220;
wire [31:0] ScanLink221;
wire [31:0] ScanLink222;
wire [31:0] ScanLink223;
wire [31:0] ScanLink224;
wire [31:0] ScanLink225;
wire [31:0] ScanLink226;
wire [31:0] ScanLink227;
wire [31:0] ScanLink228;
wire [31:0] ScanLink229;
wire [31:0] ScanLink230;
wire [31:0] ScanLink231;
wire [31:0] ScanLink232;
wire [31:0] ScanLink233;
wire [31:0] ScanLink234;
wire [31:0] ScanLink235;
wire [31:0] ScanLink236;
wire [31:0] ScanLink237;
wire [31:0] ScanLink238;
wire [31:0] ScanLink239;
wire [31:0] ScanLink240;
wire [31:0] ScanLink241;
wire [31:0] ScanLink242;
wire [31:0] ScanLink243;
wire [31:0] ScanLink244;
wire [31:0] ScanLink245;
wire [31:0] ScanLink246;
wire [31:0] ScanLink247;
wire [31:0] ScanLink248;
wire [31:0] ScanLink249;
wire [31:0] ScanLink250;
wire [31:0] ScanLink251;
wire [31:0] ScanLink252;
wire [31:0] ScanLink253;
wire [31:0] ScanLink254;
wire [31:0] ScanLink255;
wire [31:0] ScanLink256;
wire [31:0] ScanLink257;
wire [31:0] ScanLink258;
wire [31:0] ScanLink259;
wire [31:0] ScanLink260;
wire [31:0] ScanLink261;
wire [31:0] ScanLink262;
wire [31:0] ScanLink263;
wire [31:0] ScanLink264;
wire [31:0] ScanLink265;
wire [31:0] ScanLink266;
wire [31:0] ScanLink267;
wire [31:0] ScanLink268;
wire [31:0] ScanLink269;
wire [31:0] ScanLink270;
wire [31:0] ScanLink271;
wire [31:0] ScanLink272;
wire [31:0] ScanLink273;
wire [31:0] ScanLink274;
wire [31:0] ScanLink275;
wire [31:0] ScanLink276;
wire [31:0] ScanLink277;
wire [31:0] ScanLink278;
wire [31:0] ScanLink279;
wire [31:0] ScanLink280;
wire [31:0] ScanLink281;
wire [31:0] ScanLink282;
wire [31:0] ScanLink283;
wire [31:0] ScanLink284;
wire [31:0] ScanLink285;
wire [31:0] ScanLink286;
wire [31:0] ScanLink287;
wire [31:0] ScanLink288;
wire [31:0] ScanLink289;
wire [31:0] ScanLink290;
wire [31:0] ScanLink291;
wire [31:0] ScanLink292;
wire [31:0] ScanLink293;
wire [31:0] ScanLink294;
wire [31:0] ScanLink295;
wire [31:0] ScanLink296;
wire [31:0] ScanLink297;
wire [31:0] ScanLink298;
wire [31:0] ScanLink299;
wire [31:0] ScanLink300;
wire [31:0] ScanLink301;
wire [31:0] ScanLink302;
wire [31:0] ScanLink303;
wire [31:0] ScanLink304;
wire [31:0] ScanLink305;
wire [31:0] ScanLink306;
wire [31:0] ScanLink307;
wire [31:0] ScanLink308;
wire [31:0] ScanLink309;
wire [31:0] ScanLink310;
wire [31:0] ScanLink311;
wire [31:0] ScanLink312;
wire [31:0] ScanLink313;
wire [31:0] ScanLink314;
wire [31:0] ScanLink315;
wire [31:0] ScanLink316;
wire [31:0] ScanLink317;
wire [31:0] ScanLink318;
wire [31:0] ScanLink319;
wire [31:0] ScanLink320;
wire [31:0] ScanLink321;
wire [31:0] ScanLink322;
wire [31:0] ScanLink323;
wire [31:0] ScanLink324;
wire [31:0] ScanLink325;
wire [31:0] ScanLink326;
wire [31:0] ScanLink327;
wire [31:0] ScanLink328;
wire [31:0] ScanLink329;
wire [31:0] ScanLink330;
wire [31:0] ScanLink331;
wire [31:0] ScanLink332;
wire [31:0] ScanLink333;
wire [31:0] ScanLink334;
wire [31:0] ScanLink335;
wire [31:0] ScanLink336;
wire [31:0] ScanLink337;
wire [31:0] ScanLink338;
wire [31:0] ScanLink339;
wire [31:0] ScanLink340;
wire [31:0] ScanLink341;
wire [31:0] ScanLink342;
wire [31:0] ScanLink343;
wire [31:0] ScanLink344;
wire [31:0] ScanLink345;
wire [31:0] ScanLink346;
wire [31:0] ScanLink347;
wire [31:0] ScanLink348;
wire [31:0] ScanLink349;
wire [31:0] ScanLink350;
wire [31:0] ScanLink351;
wire [31:0] ScanLink352;
wire [31:0] ScanLink353;
wire [31:0] ScanLink354;
wire [31:0] ScanLink355;
wire [31:0] ScanLink356;
wire [31:0] ScanLink357;
wire [31:0] ScanLink358;
wire [31:0] ScanLink359;
wire [31:0] ScanLink360;
wire [31:0] ScanLink361;
wire [31:0] ScanLink362;
wire [31:0] ScanLink363;
wire [31:0] ScanLink364;
wire [31:0] ScanLink365;
wire [31:0] ScanLink366;
wire [31:0] ScanLink367;
wire [31:0] ScanLink368;
wire [31:0] ScanLink369;
wire [31:0] ScanLink370;
wire [31:0] ScanLink371;
wire [31:0] ScanLink372;
wire [31:0] ScanLink373;
wire [31:0] ScanLink374;
wire [31:0] ScanLink375;
wire [31:0] ScanLink376;
wire [31:0] ScanLink377;
wire [31:0] ScanLink378;
wire [31:0] ScanLink379;
wire [31:0] ScanLink380;
wire [31:0] ScanLink381;
wire [31:0] ScanLink382;
wire [31:0] ScanLink383;
wire [31:0] ScanLink384;
wire [31:0] ScanLink385;
wire [31:0] ScanLink386;
wire [31:0] ScanLink387;
wire [31:0] ScanLink388;
wire [31:0] ScanLink389;
wire [31:0] ScanLink390;
wire [31:0] ScanLink391;
wire [31:0] ScanLink392;
wire [31:0] ScanLink393;
wire [31:0] ScanLink394;
wire [31:0] ScanLink395;
wire [31:0] ScanLink396;
wire [31:0] ScanLink397;
wire [31:0] ScanLink398;
wire [31:0] ScanLink399;
wire [31:0] ScanLink400;
wire [31:0] ScanLink401;
wire [31:0] ScanLink402;
wire [31:0] ScanLink403;
wire [31:0] ScanLink404;
wire [31:0] ScanLink405;
wire [31:0] ScanLink406;
wire [31:0] ScanLink407;
wire [31:0] ScanLink408;
wire [31:0] ScanLink409;
wire [31:0] ScanLink410;
wire [31:0] ScanLink411;
wire [31:0] ScanLink412;
wire [31:0] ScanLink413;
wire [31:0] ScanLink414;
wire [31:0] ScanLink415;
wire [31:0] ScanLink416;
wire [31:0] ScanLink417;
wire [31:0] ScanLink418;
wire [31:0] ScanLink419;
wire [31:0] ScanLink420;
wire [31:0] ScanLink421;
wire [31:0] ScanLink422;
wire [31:0] ScanLink423;
wire [31:0] ScanLink424;
wire [31:0] ScanLink425;
wire [31:0] ScanLink426;
wire [31:0] ScanLink427;
wire [31:0] ScanLink428;
wire [31:0] ScanLink429;
wire [31:0] ScanLink430;
wire [31:0] ScanLink431;
wire [31:0] ScanLink432;
wire [31:0] ScanLink433;
wire [31:0] ScanLink434;
wire [31:0] ScanLink435;
wire [31:0] ScanLink436;
wire [31:0] ScanLink437;
wire [31:0] ScanLink438;
wire [31:0] ScanLink439;
wire [31:0] ScanLink440;
wire [31:0] ScanLink441;
wire [31:0] ScanLink442;
wire [31:0] ScanLink443;
wire [31:0] ScanLink444;
wire [31:0] ScanLink445;
wire [31:0] ScanLink446;
wire [31:0] ScanLink447;
wire [31:0] ScanLink448;
wire [31:0] ScanLink449;
wire [31:0] ScanLink450;
wire [31:0] ScanLink451;
wire [31:0] ScanLink452;
wire [31:0] ScanLink453;
wire [31:0] ScanLink454;
wire [31:0] ScanLink455;
wire [31:0] ScanLink456;
wire [31:0] ScanLink457;
wire [31:0] ScanLink458;
wire [31:0] ScanLink459;
wire [31:0] ScanLink460;
wire [31:0] ScanLink461;
wire [31:0] ScanLink462;
wire [31:0] ScanLink463;
wire [31:0] ScanLink464;
wire [31:0] ScanLink465;
wire [31:0] ScanLink466;
wire [31:0] ScanLink467;
wire [31:0] ScanLink468;
wire [31:0] ScanLink469;
wire [31:0] ScanLink470;
wire [31:0] ScanLink471;
wire [31:0] ScanLink472;
wire [31:0] ScanLink473;
wire [31:0] ScanLink474;
wire [31:0] ScanLink475;
wire [31:0] ScanLink476;
wire [31:0] ScanLink477;
wire [31:0] ScanLink478;
wire [31:0] ScanLink479;
wire [31:0] ScanLink480;
wire [31:0] ScanLink481;
wire [31:0] ScanLink482;
wire [31:0] ScanLink483;
wire [31:0] ScanLink484;
wire [31:0] ScanLink485;
wire [31:0] ScanLink486;
wire [31:0] ScanLink487;
wire [31:0] ScanLink488;
wire [31:0] ScanLink489;
wire [31:0] ScanLink490;
wire [31:0] ScanLink491;
wire [31:0] ScanLink492;
wire [31:0] ScanLink493;
wire [31:0] ScanLink494;
wire [31:0] ScanLink495;
wire [31:0] ScanLink496;
wire [31:0] ScanLink497;
wire [31:0] ScanLink498;
wire [31:0] ScanLink499;
wire [31:0] ScanLink500;
wire [31:0] ScanLink501;
wire [31:0] ScanLink502;
wire [31:0] ScanLink503;
wire [31:0] ScanLink504;
wire [31:0] ScanLink505;
wire [31:0] ScanLink506;
wire [31:0] ScanLink507;
wire [31:0] ScanLink508;
wire [31:0] ScanLink509;
wire [31:0] ScanLink510;
wire [31:0] ScanLink511;
wire [31:0] ScanLink512;
BubbleSort_Node #( 32 ) BSN1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn0), .BIn(wBIn0), .HiOut(wRegInA0), .LoOut(wAMid0) );
BubbleSort_Node #( 32 ) BSN1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn1), .BIn(wBIn1), .HiOut(wBMid0), .LoOut(wAMid1) );
BubbleSort_Node #( 32 ) BSN1_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn2), .BIn(wBIn2), .HiOut(wBMid1), .LoOut(wAMid2) );
BubbleSort_Node #( 32 ) BSN1_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn3), .BIn(wBIn3), .HiOut(wBMid2), .LoOut(wAMid3) );
BubbleSort_Node #( 32 ) BSN1_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn4), .BIn(wBIn4), .HiOut(wBMid3), .LoOut(wAMid4) );
BubbleSort_Node #( 32 ) BSN1_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn5), .BIn(wBIn5), .HiOut(wBMid4), .LoOut(wAMid5) );
BubbleSort_Node #( 32 ) BSN1_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn6), .BIn(wBIn6), .HiOut(wBMid5), .LoOut(wAMid6) );
BubbleSort_Node #( 32 ) BSN1_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn7), .BIn(wBIn7), .HiOut(wBMid6), .LoOut(wAMid7) );
BubbleSort_Node #( 32 ) BSN1_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn8), .BIn(wBIn8), .HiOut(wBMid7), .LoOut(wAMid8) );
BubbleSort_Node #( 32 ) BSN1_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn9), .BIn(wBIn9), .HiOut(wBMid8), .LoOut(wAMid9) );
BubbleSort_Node #( 32 ) BSN1_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn10), .BIn(wBIn10), .HiOut(wBMid9), .LoOut(wAMid10) );
BubbleSort_Node #( 32 ) BSN1_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn11), .BIn(wBIn11), .HiOut(wBMid10), .LoOut(wAMid11) );
BubbleSort_Node #( 32 ) BSN1_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn12), .BIn(wBIn12), .HiOut(wBMid11), .LoOut(wAMid12) );
BubbleSort_Node #( 32 ) BSN1_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn13), .BIn(wBIn13), .HiOut(wBMid12), .LoOut(wAMid13) );
BubbleSort_Node #( 32 ) BSN1_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn14), .BIn(wBIn14), .HiOut(wBMid13), .LoOut(wAMid14) );
BubbleSort_Node #( 32 ) BSN1_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn15), .BIn(wBIn15), .HiOut(wBMid14), .LoOut(wAMid15) );
BubbleSort_Node #( 32 ) BSN1_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn16), .BIn(wBIn16), .HiOut(wBMid15), .LoOut(wAMid16) );
BubbleSort_Node #( 32 ) BSN1_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn17), .BIn(wBIn17), .HiOut(wBMid16), .LoOut(wAMid17) );
BubbleSort_Node #( 32 ) BSN1_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn18), .BIn(wBIn18), .HiOut(wBMid17), .LoOut(wAMid18) );
BubbleSort_Node #( 32 ) BSN1_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn19), .BIn(wBIn19), .HiOut(wBMid18), .LoOut(wAMid19) );
BubbleSort_Node #( 32 ) BSN1_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn20), .BIn(wBIn20), .HiOut(wBMid19), .LoOut(wAMid20) );
BubbleSort_Node #( 32 ) BSN1_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn21), .BIn(wBIn21), .HiOut(wBMid20), .LoOut(wAMid21) );
BubbleSort_Node #( 32 ) BSN1_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn22), .BIn(wBIn22), .HiOut(wBMid21), .LoOut(wAMid22) );
BubbleSort_Node #( 32 ) BSN1_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn23), .BIn(wBIn23), .HiOut(wBMid22), .LoOut(wAMid23) );
BubbleSort_Node #( 32 ) BSN1_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn24), .BIn(wBIn24), .HiOut(wBMid23), .LoOut(wAMid24) );
BubbleSort_Node #( 32 ) BSN1_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn25), .BIn(wBIn25), .HiOut(wBMid24), .LoOut(wAMid25) );
BubbleSort_Node #( 32 ) BSN1_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn26), .BIn(wBIn26), .HiOut(wBMid25), .LoOut(wAMid26) );
BubbleSort_Node #( 32 ) BSN1_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn27), .BIn(wBIn27), .HiOut(wBMid26), .LoOut(wAMid27) );
BubbleSort_Node #( 32 ) BSN1_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn28), .BIn(wBIn28), .HiOut(wBMid27), .LoOut(wAMid28) );
BubbleSort_Node #( 32 ) BSN1_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn29), .BIn(wBIn29), .HiOut(wBMid28), .LoOut(wAMid29) );
BubbleSort_Node #( 32 ) BSN1_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn30), .BIn(wBIn30), .HiOut(wBMid29), .LoOut(wAMid30) );
BubbleSort_Node #( 32 ) BSN1_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn31), .BIn(wBIn31), .HiOut(wBMid30), .LoOut(wAMid31) );
BubbleSort_Node #( 32 ) BSN1_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn32), .BIn(wBIn32), .HiOut(wBMid31), .LoOut(wAMid32) );
BubbleSort_Node #( 32 ) BSN1_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn33), .BIn(wBIn33), .HiOut(wBMid32), .LoOut(wAMid33) );
BubbleSort_Node #( 32 ) BSN1_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn34), .BIn(wBIn34), .HiOut(wBMid33), .LoOut(wAMid34) );
BubbleSort_Node #( 32 ) BSN1_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn35), .BIn(wBIn35), .HiOut(wBMid34), .LoOut(wAMid35) );
BubbleSort_Node #( 32 ) BSN1_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn36), .BIn(wBIn36), .HiOut(wBMid35), .LoOut(wAMid36) );
BubbleSort_Node #( 32 ) BSN1_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn37), .BIn(wBIn37), .HiOut(wBMid36), .LoOut(wAMid37) );
BubbleSort_Node #( 32 ) BSN1_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn38), .BIn(wBIn38), .HiOut(wBMid37), .LoOut(wAMid38) );
BubbleSort_Node #( 32 ) BSN1_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn39), .BIn(wBIn39), .HiOut(wBMid38), .LoOut(wAMid39) );
BubbleSort_Node #( 32 ) BSN1_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn40), .BIn(wBIn40), .HiOut(wBMid39), .LoOut(wAMid40) );
BubbleSort_Node #( 32 ) BSN1_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn41), .BIn(wBIn41), .HiOut(wBMid40), .LoOut(wAMid41) );
BubbleSort_Node #( 32 ) BSN1_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn42), .BIn(wBIn42), .HiOut(wBMid41), .LoOut(wAMid42) );
BubbleSort_Node #( 32 ) BSN1_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn43), .BIn(wBIn43), .HiOut(wBMid42), .LoOut(wAMid43) );
BubbleSort_Node #( 32 ) BSN1_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn44), .BIn(wBIn44), .HiOut(wBMid43), .LoOut(wAMid44) );
BubbleSort_Node #( 32 ) BSN1_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn45), .BIn(wBIn45), .HiOut(wBMid44), .LoOut(wAMid45) );
BubbleSort_Node #( 32 ) BSN1_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn46), .BIn(wBIn46), .HiOut(wBMid45), .LoOut(wAMid46) );
BubbleSort_Node #( 32 ) BSN1_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn47), .BIn(wBIn47), .HiOut(wBMid46), .LoOut(wAMid47) );
BubbleSort_Node #( 32 ) BSN1_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn48), .BIn(wBIn48), .HiOut(wBMid47), .LoOut(wAMid48) );
BubbleSort_Node #( 32 ) BSN1_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn49), .BIn(wBIn49), .HiOut(wBMid48), .LoOut(wAMid49) );
BubbleSort_Node #( 32 ) BSN1_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn50), .BIn(wBIn50), .HiOut(wBMid49), .LoOut(wAMid50) );
BubbleSort_Node #( 32 ) BSN1_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn51), .BIn(wBIn51), .HiOut(wBMid50), .LoOut(wAMid51) );
BubbleSort_Node #( 32 ) BSN1_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn52), .BIn(wBIn52), .HiOut(wBMid51), .LoOut(wAMid52) );
BubbleSort_Node #( 32 ) BSN1_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn53), .BIn(wBIn53), .HiOut(wBMid52), .LoOut(wAMid53) );
BubbleSort_Node #( 32 ) BSN1_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn54), .BIn(wBIn54), .HiOut(wBMid53), .LoOut(wAMid54) );
BubbleSort_Node #( 32 ) BSN1_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn55), .BIn(wBIn55), .HiOut(wBMid54), .LoOut(wAMid55) );
BubbleSort_Node #( 32 ) BSN1_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn56), .BIn(wBIn56), .HiOut(wBMid55), .LoOut(wAMid56) );
BubbleSort_Node #( 32 ) BSN1_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn57), .BIn(wBIn57), .HiOut(wBMid56), .LoOut(wAMid57) );
BubbleSort_Node #( 32 ) BSN1_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn58), .BIn(wBIn58), .HiOut(wBMid57), .LoOut(wAMid58) );
BubbleSort_Node #( 32 ) BSN1_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn59), .BIn(wBIn59), .HiOut(wBMid58), .LoOut(wAMid59) );
BubbleSort_Node #( 32 ) BSN1_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn60), .BIn(wBIn60), .HiOut(wBMid59), .LoOut(wAMid60) );
BubbleSort_Node #( 32 ) BSN1_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn61), .BIn(wBIn61), .HiOut(wBMid60), .LoOut(wAMid61) );
BubbleSort_Node #( 32 ) BSN1_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn62), .BIn(wBIn62), .HiOut(wBMid61), .LoOut(wAMid62) );
BubbleSort_Node #( 32 ) BSN1_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn63), .BIn(wBIn63), .HiOut(wBMid62), .LoOut(wAMid63) );
BubbleSort_Node #( 32 ) BSN1_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn64), .BIn(wBIn64), .HiOut(wBMid63), .LoOut(wAMid64) );
BubbleSort_Node #( 32 ) BSN1_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn65), .BIn(wBIn65), .HiOut(wBMid64), .LoOut(wAMid65) );
BubbleSort_Node #( 32 ) BSN1_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn66), .BIn(wBIn66), .HiOut(wBMid65), .LoOut(wAMid66) );
BubbleSort_Node #( 32 ) BSN1_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn67), .BIn(wBIn67), .HiOut(wBMid66), .LoOut(wAMid67) );
BubbleSort_Node #( 32 ) BSN1_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn68), .BIn(wBIn68), .HiOut(wBMid67), .LoOut(wAMid68) );
BubbleSort_Node #( 32 ) BSN1_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn69), .BIn(wBIn69), .HiOut(wBMid68), .LoOut(wAMid69) );
BubbleSort_Node #( 32 ) BSN1_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn70), .BIn(wBIn70), .HiOut(wBMid69), .LoOut(wAMid70) );
BubbleSort_Node #( 32 ) BSN1_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn71), .BIn(wBIn71), .HiOut(wBMid70), .LoOut(wAMid71) );
BubbleSort_Node #( 32 ) BSN1_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn72), .BIn(wBIn72), .HiOut(wBMid71), .LoOut(wAMid72) );
BubbleSort_Node #( 32 ) BSN1_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn73), .BIn(wBIn73), .HiOut(wBMid72), .LoOut(wAMid73) );
BubbleSort_Node #( 32 ) BSN1_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn74), .BIn(wBIn74), .HiOut(wBMid73), .LoOut(wAMid74) );
BubbleSort_Node #( 32 ) BSN1_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn75), .BIn(wBIn75), .HiOut(wBMid74), .LoOut(wAMid75) );
BubbleSort_Node #( 32 ) BSN1_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn76), .BIn(wBIn76), .HiOut(wBMid75), .LoOut(wAMid76) );
BubbleSort_Node #( 32 ) BSN1_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn77), .BIn(wBIn77), .HiOut(wBMid76), .LoOut(wAMid77) );
BubbleSort_Node #( 32 ) BSN1_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn78), .BIn(wBIn78), .HiOut(wBMid77), .LoOut(wAMid78) );
BubbleSort_Node #( 32 ) BSN1_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn79), .BIn(wBIn79), .HiOut(wBMid78), .LoOut(wAMid79) );
BubbleSort_Node #( 32 ) BSN1_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn80), .BIn(wBIn80), .HiOut(wBMid79), .LoOut(wAMid80) );
BubbleSort_Node #( 32 ) BSN1_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn81), .BIn(wBIn81), .HiOut(wBMid80), .LoOut(wAMid81) );
BubbleSort_Node #( 32 ) BSN1_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn82), .BIn(wBIn82), .HiOut(wBMid81), .LoOut(wAMid82) );
BubbleSort_Node #( 32 ) BSN1_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn83), .BIn(wBIn83), .HiOut(wBMid82), .LoOut(wAMid83) );
BubbleSort_Node #( 32 ) BSN1_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn84), .BIn(wBIn84), .HiOut(wBMid83), .LoOut(wAMid84) );
BubbleSort_Node #( 32 ) BSN1_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn85), .BIn(wBIn85), .HiOut(wBMid84), .LoOut(wAMid85) );
BubbleSort_Node #( 32 ) BSN1_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn86), .BIn(wBIn86), .HiOut(wBMid85), .LoOut(wAMid86) );
BubbleSort_Node #( 32 ) BSN1_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn87), .BIn(wBIn87), .HiOut(wBMid86), .LoOut(wAMid87) );
BubbleSort_Node #( 32 ) BSN1_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn88), .BIn(wBIn88), .HiOut(wBMid87), .LoOut(wAMid88) );
BubbleSort_Node #( 32 ) BSN1_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn89), .BIn(wBIn89), .HiOut(wBMid88), .LoOut(wAMid89) );
BubbleSort_Node #( 32 ) BSN1_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn90), .BIn(wBIn90), .HiOut(wBMid89), .LoOut(wAMid90) );
BubbleSort_Node #( 32 ) BSN1_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn91), .BIn(wBIn91), .HiOut(wBMid90), .LoOut(wAMid91) );
BubbleSort_Node #( 32 ) BSN1_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn92), .BIn(wBIn92), .HiOut(wBMid91), .LoOut(wAMid92) );
BubbleSort_Node #( 32 ) BSN1_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn93), .BIn(wBIn93), .HiOut(wBMid92), .LoOut(wAMid93) );
BubbleSort_Node #( 32 ) BSN1_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn94), .BIn(wBIn94), .HiOut(wBMid93), .LoOut(wAMid94) );
BubbleSort_Node #( 32 ) BSN1_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn95), .BIn(wBIn95), .HiOut(wBMid94), .LoOut(wAMid95) );
BubbleSort_Node #( 32 ) BSN1_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn96), .BIn(wBIn96), .HiOut(wBMid95), .LoOut(wAMid96) );
BubbleSort_Node #( 32 ) BSN1_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn97), .BIn(wBIn97), .HiOut(wBMid96), .LoOut(wAMid97) );
BubbleSort_Node #( 32 ) BSN1_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn98), .BIn(wBIn98), .HiOut(wBMid97), .LoOut(wAMid98) );
BubbleSort_Node #( 32 ) BSN1_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn99), .BIn(wBIn99), .HiOut(wBMid98), .LoOut(wAMid99) );
BubbleSort_Node #( 32 ) BSN1_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn100), .BIn(wBIn100), .HiOut(wBMid99), .LoOut(wAMid100) );
BubbleSort_Node #( 32 ) BSN1_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn101), .BIn(wBIn101), .HiOut(wBMid100), .LoOut(wAMid101) );
BubbleSort_Node #( 32 ) BSN1_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn102), .BIn(wBIn102), .HiOut(wBMid101), .LoOut(wAMid102) );
BubbleSort_Node #( 32 ) BSN1_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn103), .BIn(wBIn103), .HiOut(wBMid102), .LoOut(wAMid103) );
BubbleSort_Node #( 32 ) BSN1_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn104), .BIn(wBIn104), .HiOut(wBMid103), .LoOut(wAMid104) );
BubbleSort_Node #( 32 ) BSN1_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn105), .BIn(wBIn105), .HiOut(wBMid104), .LoOut(wAMid105) );
BubbleSort_Node #( 32 ) BSN1_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn106), .BIn(wBIn106), .HiOut(wBMid105), .LoOut(wAMid106) );
BubbleSort_Node #( 32 ) BSN1_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn107), .BIn(wBIn107), .HiOut(wBMid106), .LoOut(wAMid107) );
BubbleSort_Node #( 32 ) BSN1_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn108), .BIn(wBIn108), .HiOut(wBMid107), .LoOut(wAMid108) );
BubbleSort_Node #( 32 ) BSN1_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn109), .BIn(wBIn109), .HiOut(wBMid108), .LoOut(wAMid109) );
BubbleSort_Node #( 32 ) BSN1_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn110), .BIn(wBIn110), .HiOut(wBMid109), .LoOut(wAMid110) );
BubbleSort_Node #( 32 ) BSN1_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn111), .BIn(wBIn111), .HiOut(wBMid110), .LoOut(wAMid111) );
BubbleSort_Node #( 32 ) BSN1_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn112), .BIn(wBIn112), .HiOut(wBMid111), .LoOut(wAMid112) );
BubbleSort_Node #( 32 ) BSN1_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn113), .BIn(wBIn113), .HiOut(wBMid112), .LoOut(wAMid113) );
BubbleSort_Node #( 32 ) BSN1_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn114), .BIn(wBIn114), .HiOut(wBMid113), .LoOut(wAMid114) );
BubbleSort_Node #( 32 ) BSN1_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn115), .BIn(wBIn115), .HiOut(wBMid114), .LoOut(wAMid115) );
BubbleSort_Node #( 32 ) BSN1_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn116), .BIn(wBIn116), .HiOut(wBMid115), .LoOut(wAMid116) );
BubbleSort_Node #( 32 ) BSN1_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn117), .BIn(wBIn117), .HiOut(wBMid116), .LoOut(wAMid117) );
BubbleSort_Node #( 32 ) BSN1_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn118), .BIn(wBIn118), .HiOut(wBMid117), .LoOut(wAMid118) );
BubbleSort_Node #( 32 ) BSN1_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn119), .BIn(wBIn119), .HiOut(wBMid118), .LoOut(wAMid119) );
BubbleSort_Node #( 32 ) BSN1_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn120), .BIn(wBIn120), .HiOut(wBMid119), .LoOut(wAMid120) );
BubbleSort_Node #( 32 ) BSN1_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn121), .BIn(wBIn121), .HiOut(wBMid120), .LoOut(wAMid121) );
BubbleSort_Node #( 32 ) BSN1_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn122), .BIn(wBIn122), .HiOut(wBMid121), .LoOut(wAMid122) );
BubbleSort_Node #( 32 ) BSN1_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn123), .BIn(wBIn123), .HiOut(wBMid122), .LoOut(wAMid123) );
BubbleSort_Node #( 32 ) BSN1_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn124), .BIn(wBIn124), .HiOut(wBMid123), .LoOut(wAMid124) );
BubbleSort_Node #( 32 ) BSN1_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn125), .BIn(wBIn125), .HiOut(wBMid124), .LoOut(wAMid125) );
BubbleSort_Node #( 32 ) BSN1_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn126), .BIn(wBIn126), .HiOut(wBMid125), .LoOut(wAMid126) );
BubbleSort_Node #( 32 ) BSN1_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn127), .BIn(wBIn127), .HiOut(wBMid126), .LoOut(wAMid127) );
BubbleSort_Node #( 32 ) BSN1_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn128), .BIn(wBIn128), .HiOut(wBMid127), .LoOut(wAMid128) );
BubbleSort_Node #( 32 ) BSN1_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn129), .BIn(wBIn129), .HiOut(wBMid128), .LoOut(wAMid129) );
BubbleSort_Node #( 32 ) BSN1_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn130), .BIn(wBIn130), .HiOut(wBMid129), .LoOut(wAMid130) );
BubbleSort_Node #( 32 ) BSN1_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn131), .BIn(wBIn131), .HiOut(wBMid130), .LoOut(wAMid131) );
BubbleSort_Node #( 32 ) BSN1_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn132), .BIn(wBIn132), .HiOut(wBMid131), .LoOut(wAMid132) );
BubbleSort_Node #( 32 ) BSN1_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn133), .BIn(wBIn133), .HiOut(wBMid132), .LoOut(wAMid133) );
BubbleSort_Node #( 32 ) BSN1_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn134), .BIn(wBIn134), .HiOut(wBMid133), .LoOut(wAMid134) );
BubbleSort_Node #( 32 ) BSN1_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn135), .BIn(wBIn135), .HiOut(wBMid134), .LoOut(wAMid135) );
BubbleSort_Node #( 32 ) BSN1_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn136), .BIn(wBIn136), .HiOut(wBMid135), .LoOut(wAMid136) );
BubbleSort_Node #( 32 ) BSN1_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn137), .BIn(wBIn137), .HiOut(wBMid136), .LoOut(wAMid137) );
BubbleSort_Node #( 32 ) BSN1_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn138), .BIn(wBIn138), .HiOut(wBMid137), .LoOut(wAMid138) );
BubbleSort_Node #( 32 ) BSN1_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn139), .BIn(wBIn139), .HiOut(wBMid138), .LoOut(wAMid139) );
BubbleSort_Node #( 32 ) BSN1_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn140), .BIn(wBIn140), .HiOut(wBMid139), .LoOut(wAMid140) );
BubbleSort_Node #( 32 ) BSN1_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn141), .BIn(wBIn141), .HiOut(wBMid140), .LoOut(wAMid141) );
BubbleSort_Node #( 32 ) BSN1_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn142), .BIn(wBIn142), .HiOut(wBMid141), .LoOut(wAMid142) );
BubbleSort_Node #( 32 ) BSN1_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn143), .BIn(wBIn143), .HiOut(wBMid142), .LoOut(wAMid143) );
BubbleSort_Node #( 32 ) BSN1_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn144), .BIn(wBIn144), .HiOut(wBMid143), .LoOut(wAMid144) );
BubbleSort_Node #( 32 ) BSN1_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn145), .BIn(wBIn145), .HiOut(wBMid144), .LoOut(wAMid145) );
BubbleSort_Node #( 32 ) BSN1_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn146), .BIn(wBIn146), .HiOut(wBMid145), .LoOut(wAMid146) );
BubbleSort_Node #( 32 ) BSN1_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn147), .BIn(wBIn147), .HiOut(wBMid146), .LoOut(wAMid147) );
BubbleSort_Node #( 32 ) BSN1_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn148), .BIn(wBIn148), .HiOut(wBMid147), .LoOut(wAMid148) );
BubbleSort_Node #( 32 ) BSN1_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn149), .BIn(wBIn149), .HiOut(wBMid148), .LoOut(wAMid149) );
BubbleSort_Node #( 32 ) BSN1_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn150), .BIn(wBIn150), .HiOut(wBMid149), .LoOut(wAMid150) );
BubbleSort_Node #( 32 ) BSN1_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn151), .BIn(wBIn151), .HiOut(wBMid150), .LoOut(wAMid151) );
BubbleSort_Node #( 32 ) BSN1_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn152), .BIn(wBIn152), .HiOut(wBMid151), .LoOut(wAMid152) );
BubbleSort_Node #( 32 ) BSN1_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn153), .BIn(wBIn153), .HiOut(wBMid152), .LoOut(wAMid153) );
BubbleSort_Node #( 32 ) BSN1_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn154), .BIn(wBIn154), .HiOut(wBMid153), .LoOut(wAMid154) );
BubbleSort_Node #( 32 ) BSN1_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn155), .BIn(wBIn155), .HiOut(wBMid154), .LoOut(wAMid155) );
BubbleSort_Node #( 32 ) BSN1_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn156), .BIn(wBIn156), .HiOut(wBMid155), .LoOut(wAMid156) );
BubbleSort_Node #( 32 ) BSN1_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn157), .BIn(wBIn157), .HiOut(wBMid156), .LoOut(wAMid157) );
BubbleSort_Node #( 32 ) BSN1_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn158), .BIn(wBIn158), .HiOut(wBMid157), .LoOut(wAMid158) );
BubbleSort_Node #( 32 ) BSN1_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn159), .BIn(wBIn159), .HiOut(wBMid158), .LoOut(wAMid159) );
BubbleSort_Node #( 32 ) BSN1_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn160), .BIn(wBIn160), .HiOut(wBMid159), .LoOut(wAMid160) );
BubbleSort_Node #( 32 ) BSN1_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn161), .BIn(wBIn161), .HiOut(wBMid160), .LoOut(wAMid161) );
BubbleSort_Node #( 32 ) BSN1_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn162), .BIn(wBIn162), .HiOut(wBMid161), .LoOut(wAMid162) );
BubbleSort_Node #( 32 ) BSN1_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn163), .BIn(wBIn163), .HiOut(wBMid162), .LoOut(wAMid163) );
BubbleSort_Node #( 32 ) BSN1_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn164), .BIn(wBIn164), .HiOut(wBMid163), .LoOut(wAMid164) );
BubbleSort_Node #( 32 ) BSN1_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn165), .BIn(wBIn165), .HiOut(wBMid164), .LoOut(wAMid165) );
BubbleSort_Node #( 32 ) BSN1_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn166), .BIn(wBIn166), .HiOut(wBMid165), .LoOut(wAMid166) );
BubbleSort_Node #( 32 ) BSN1_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn167), .BIn(wBIn167), .HiOut(wBMid166), .LoOut(wAMid167) );
BubbleSort_Node #( 32 ) BSN1_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn168), .BIn(wBIn168), .HiOut(wBMid167), .LoOut(wAMid168) );
BubbleSort_Node #( 32 ) BSN1_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn169), .BIn(wBIn169), .HiOut(wBMid168), .LoOut(wAMid169) );
BubbleSort_Node #( 32 ) BSN1_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn170), .BIn(wBIn170), .HiOut(wBMid169), .LoOut(wAMid170) );
BubbleSort_Node #( 32 ) BSN1_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn171), .BIn(wBIn171), .HiOut(wBMid170), .LoOut(wAMid171) );
BubbleSort_Node #( 32 ) BSN1_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn172), .BIn(wBIn172), .HiOut(wBMid171), .LoOut(wAMid172) );
BubbleSort_Node #( 32 ) BSN1_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn173), .BIn(wBIn173), .HiOut(wBMid172), .LoOut(wAMid173) );
BubbleSort_Node #( 32 ) BSN1_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn174), .BIn(wBIn174), .HiOut(wBMid173), .LoOut(wAMid174) );
BubbleSort_Node #( 32 ) BSN1_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn175), .BIn(wBIn175), .HiOut(wBMid174), .LoOut(wAMid175) );
BubbleSort_Node #( 32 ) BSN1_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn176), .BIn(wBIn176), .HiOut(wBMid175), .LoOut(wAMid176) );
BubbleSort_Node #( 32 ) BSN1_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn177), .BIn(wBIn177), .HiOut(wBMid176), .LoOut(wAMid177) );
BubbleSort_Node #( 32 ) BSN1_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn178), .BIn(wBIn178), .HiOut(wBMid177), .LoOut(wAMid178) );
BubbleSort_Node #( 32 ) BSN1_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn179), .BIn(wBIn179), .HiOut(wBMid178), .LoOut(wAMid179) );
BubbleSort_Node #( 32 ) BSN1_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn180), .BIn(wBIn180), .HiOut(wBMid179), .LoOut(wAMid180) );
BubbleSort_Node #( 32 ) BSN1_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn181), .BIn(wBIn181), .HiOut(wBMid180), .LoOut(wAMid181) );
BubbleSort_Node #( 32 ) BSN1_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn182), .BIn(wBIn182), .HiOut(wBMid181), .LoOut(wAMid182) );
BubbleSort_Node #( 32 ) BSN1_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn183), .BIn(wBIn183), .HiOut(wBMid182), .LoOut(wAMid183) );
BubbleSort_Node #( 32 ) BSN1_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn184), .BIn(wBIn184), .HiOut(wBMid183), .LoOut(wAMid184) );
BubbleSort_Node #( 32 ) BSN1_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn185), .BIn(wBIn185), .HiOut(wBMid184), .LoOut(wAMid185) );
BubbleSort_Node #( 32 ) BSN1_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn186), .BIn(wBIn186), .HiOut(wBMid185), .LoOut(wAMid186) );
BubbleSort_Node #( 32 ) BSN1_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn187), .BIn(wBIn187), .HiOut(wBMid186), .LoOut(wAMid187) );
BubbleSort_Node #( 32 ) BSN1_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn188), .BIn(wBIn188), .HiOut(wBMid187), .LoOut(wAMid188) );
BubbleSort_Node #( 32 ) BSN1_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn189), .BIn(wBIn189), .HiOut(wBMid188), .LoOut(wAMid189) );
BubbleSort_Node #( 32 ) BSN1_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn190), .BIn(wBIn190), .HiOut(wBMid189), .LoOut(wAMid190) );
BubbleSort_Node #( 32 ) BSN1_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn191), .BIn(wBIn191), .HiOut(wBMid190), .LoOut(wAMid191) );
BubbleSort_Node #( 32 ) BSN1_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn192), .BIn(wBIn192), .HiOut(wBMid191), .LoOut(wAMid192) );
BubbleSort_Node #( 32 ) BSN1_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn193), .BIn(wBIn193), .HiOut(wBMid192), .LoOut(wAMid193) );
BubbleSort_Node #( 32 ) BSN1_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn194), .BIn(wBIn194), .HiOut(wBMid193), .LoOut(wAMid194) );
BubbleSort_Node #( 32 ) BSN1_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn195), .BIn(wBIn195), .HiOut(wBMid194), .LoOut(wAMid195) );
BubbleSort_Node #( 32 ) BSN1_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn196), .BIn(wBIn196), .HiOut(wBMid195), .LoOut(wAMid196) );
BubbleSort_Node #( 32 ) BSN1_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn197), .BIn(wBIn197), .HiOut(wBMid196), .LoOut(wAMid197) );
BubbleSort_Node #( 32 ) BSN1_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn198), .BIn(wBIn198), .HiOut(wBMid197), .LoOut(wAMid198) );
BubbleSort_Node #( 32 ) BSN1_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn199), .BIn(wBIn199), .HiOut(wBMid198), .LoOut(wAMid199) );
BubbleSort_Node #( 32 ) BSN1_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn200), .BIn(wBIn200), .HiOut(wBMid199), .LoOut(wAMid200) );
BubbleSort_Node #( 32 ) BSN1_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn201), .BIn(wBIn201), .HiOut(wBMid200), .LoOut(wAMid201) );
BubbleSort_Node #( 32 ) BSN1_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn202), .BIn(wBIn202), .HiOut(wBMid201), .LoOut(wAMid202) );
BubbleSort_Node #( 32 ) BSN1_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn203), .BIn(wBIn203), .HiOut(wBMid202), .LoOut(wAMid203) );
BubbleSort_Node #( 32 ) BSN1_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn204), .BIn(wBIn204), .HiOut(wBMid203), .LoOut(wAMid204) );
BubbleSort_Node #( 32 ) BSN1_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn205), .BIn(wBIn205), .HiOut(wBMid204), .LoOut(wAMid205) );
BubbleSort_Node #( 32 ) BSN1_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn206), .BIn(wBIn206), .HiOut(wBMid205), .LoOut(wAMid206) );
BubbleSort_Node #( 32 ) BSN1_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn207), .BIn(wBIn207), .HiOut(wBMid206), .LoOut(wAMid207) );
BubbleSort_Node #( 32 ) BSN1_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn208), .BIn(wBIn208), .HiOut(wBMid207), .LoOut(wAMid208) );
BubbleSort_Node #( 32 ) BSN1_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn209), .BIn(wBIn209), .HiOut(wBMid208), .LoOut(wAMid209) );
BubbleSort_Node #( 32 ) BSN1_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn210), .BIn(wBIn210), .HiOut(wBMid209), .LoOut(wAMid210) );
BubbleSort_Node #( 32 ) BSN1_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn211), .BIn(wBIn211), .HiOut(wBMid210), .LoOut(wAMid211) );
BubbleSort_Node #( 32 ) BSN1_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn212), .BIn(wBIn212), .HiOut(wBMid211), .LoOut(wAMid212) );
BubbleSort_Node #( 32 ) BSN1_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn213), .BIn(wBIn213), .HiOut(wBMid212), .LoOut(wAMid213) );
BubbleSort_Node #( 32 ) BSN1_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn214), .BIn(wBIn214), .HiOut(wBMid213), .LoOut(wAMid214) );
BubbleSort_Node #( 32 ) BSN1_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn215), .BIn(wBIn215), .HiOut(wBMid214), .LoOut(wAMid215) );
BubbleSort_Node #( 32 ) BSN1_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn216), .BIn(wBIn216), .HiOut(wBMid215), .LoOut(wAMid216) );
BubbleSort_Node #( 32 ) BSN1_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn217), .BIn(wBIn217), .HiOut(wBMid216), .LoOut(wAMid217) );
BubbleSort_Node #( 32 ) BSN1_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn218), .BIn(wBIn218), .HiOut(wBMid217), .LoOut(wAMid218) );
BubbleSort_Node #( 32 ) BSN1_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn219), .BIn(wBIn219), .HiOut(wBMid218), .LoOut(wAMid219) );
BubbleSort_Node #( 32 ) BSN1_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn220), .BIn(wBIn220), .HiOut(wBMid219), .LoOut(wAMid220) );
BubbleSort_Node #( 32 ) BSN1_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn221), .BIn(wBIn221), .HiOut(wBMid220), .LoOut(wAMid221) );
BubbleSort_Node #( 32 ) BSN1_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn222), .BIn(wBIn222), .HiOut(wBMid221), .LoOut(wAMid222) );
BubbleSort_Node #( 32 ) BSN1_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn223), .BIn(wBIn223), .HiOut(wBMid222), .LoOut(wAMid223) );
BubbleSort_Node #( 32 ) BSN1_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn224), .BIn(wBIn224), .HiOut(wBMid223), .LoOut(wAMid224) );
BubbleSort_Node #( 32 ) BSN1_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn225), .BIn(wBIn225), .HiOut(wBMid224), .LoOut(wAMid225) );
BubbleSort_Node #( 32 ) BSN1_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn226), .BIn(wBIn226), .HiOut(wBMid225), .LoOut(wAMid226) );
BubbleSort_Node #( 32 ) BSN1_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn227), .BIn(wBIn227), .HiOut(wBMid226), .LoOut(wAMid227) );
BubbleSort_Node #( 32 ) BSN1_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn228), .BIn(wBIn228), .HiOut(wBMid227), .LoOut(wAMid228) );
BubbleSort_Node #( 32 ) BSN1_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn229), .BIn(wBIn229), .HiOut(wBMid228), .LoOut(wAMid229) );
BubbleSort_Node #( 32 ) BSN1_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn230), .BIn(wBIn230), .HiOut(wBMid229), .LoOut(wAMid230) );
BubbleSort_Node #( 32 ) BSN1_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn231), .BIn(wBIn231), .HiOut(wBMid230), .LoOut(wAMid231) );
BubbleSort_Node #( 32 ) BSN1_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn232), .BIn(wBIn232), .HiOut(wBMid231), .LoOut(wAMid232) );
BubbleSort_Node #( 32 ) BSN1_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn233), .BIn(wBIn233), .HiOut(wBMid232), .LoOut(wAMid233) );
BubbleSort_Node #( 32 ) BSN1_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn234), .BIn(wBIn234), .HiOut(wBMid233), .LoOut(wAMid234) );
BubbleSort_Node #( 32 ) BSN1_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn235), .BIn(wBIn235), .HiOut(wBMid234), .LoOut(wAMid235) );
BubbleSort_Node #( 32 ) BSN1_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn236), .BIn(wBIn236), .HiOut(wBMid235), .LoOut(wAMid236) );
BubbleSort_Node #( 32 ) BSN1_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn237), .BIn(wBIn237), .HiOut(wBMid236), .LoOut(wAMid237) );
BubbleSort_Node #( 32 ) BSN1_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn238), .BIn(wBIn238), .HiOut(wBMid237), .LoOut(wAMid238) );
BubbleSort_Node #( 32 ) BSN1_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn239), .BIn(wBIn239), .HiOut(wBMid238), .LoOut(wAMid239) );
BubbleSort_Node #( 32 ) BSN1_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn240), .BIn(wBIn240), .HiOut(wBMid239), .LoOut(wAMid240) );
BubbleSort_Node #( 32 ) BSN1_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn241), .BIn(wBIn241), .HiOut(wBMid240), .LoOut(wAMid241) );
BubbleSort_Node #( 32 ) BSN1_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn242), .BIn(wBIn242), .HiOut(wBMid241), .LoOut(wAMid242) );
BubbleSort_Node #( 32 ) BSN1_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn243), .BIn(wBIn243), .HiOut(wBMid242), .LoOut(wAMid243) );
BubbleSort_Node #( 32 ) BSN1_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn244), .BIn(wBIn244), .HiOut(wBMid243), .LoOut(wAMid244) );
BubbleSort_Node #( 32 ) BSN1_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn245), .BIn(wBIn245), .HiOut(wBMid244), .LoOut(wAMid245) );
BubbleSort_Node #( 32 ) BSN1_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn246), .BIn(wBIn246), .HiOut(wBMid245), .LoOut(wAMid246) );
BubbleSort_Node #( 32 ) BSN1_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn247), .BIn(wBIn247), .HiOut(wBMid246), .LoOut(wAMid247) );
BubbleSort_Node #( 32 ) BSN1_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn248), .BIn(wBIn248), .HiOut(wBMid247), .LoOut(wAMid248) );
BubbleSort_Node #( 32 ) BSN1_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn249), .BIn(wBIn249), .HiOut(wBMid248), .LoOut(wAMid249) );
BubbleSort_Node #( 32 ) BSN1_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn250), .BIn(wBIn250), .HiOut(wBMid249), .LoOut(wAMid250) );
BubbleSort_Node #( 32 ) BSN1_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn251), .BIn(wBIn251), .HiOut(wBMid250), .LoOut(wAMid251) );
BubbleSort_Node #( 32 ) BSN1_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn252), .BIn(wBIn252), .HiOut(wBMid251), .LoOut(wAMid252) );
BubbleSort_Node #( 32 ) BSN1_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn253), .BIn(wBIn253), .HiOut(wBMid252), .LoOut(wAMid253) );
BubbleSort_Node #( 32 ) BSN1_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn254), .BIn(wBIn254), .HiOut(wBMid253), .LoOut(wAMid254) );
BubbleSort_Node #( 32 ) BSN1_255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAIn255), .BIn(wBIn255), .HiOut(wBMid254), .LoOut(wRegInB255) );
BubbleSort_Node #( 32 ) BSN2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid0), .BIn(wBMid0), .HiOut(wRegInB0), .LoOut(wRegInA1) );
BubbleSort_Node #( 32 ) BSN2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid1), .BIn(wBMid1), .HiOut(wRegInB1), .LoOut(wRegInA2) );
BubbleSort_Node #( 32 ) BSN2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid2), .BIn(wBMid2), .HiOut(wRegInB2), .LoOut(wRegInA3) );
BubbleSort_Node #( 32 ) BSN2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid3), .BIn(wBMid3), .HiOut(wRegInB3), .LoOut(wRegInA4) );
BubbleSort_Node #( 32 ) BSN2_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid4), .BIn(wBMid4), .HiOut(wRegInB4), .LoOut(wRegInA5) );
BubbleSort_Node #( 32 ) BSN2_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid5), .BIn(wBMid5), .HiOut(wRegInB5), .LoOut(wRegInA6) );
BubbleSort_Node #( 32 ) BSN2_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid6), .BIn(wBMid6), .HiOut(wRegInB6), .LoOut(wRegInA7) );
BubbleSort_Node #( 32 ) BSN2_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid7), .BIn(wBMid7), .HiOut(wRegInB7), .LoOut(wRegInA8) );
BubbleSort_Node #( 32 ) BSN2_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid8), .BIn(wBMid8), .HiOut(wRegInB8), .LoOut(wRegInA9) );
BubbleSort_Node #( 32 ) BSN2_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid9), .BIn(wBMid9), .HiOut(wRegInB9), .LoOut(wRegInA10) );
BubbleSort_Node #( 32 ) BSN2_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid10), .BIn(wBMid10), .HiOut(wRegInB10), .LoOut(wRegInA11) );
BubbleSort_Node #( 32 ) BSN2_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid11), .BIn(wBMid11), .HiOut(wRegInB11), .LoOut(wRegInA12) );
BubbleSort_Node #( 32 ) BSN2_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid12), .BIn(wBMid12), .HiOut(wRegInB12), .LoOut(wRegInA13) );
BubbleSort_Node #( 32 ) BSN2_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid13), .BIn(wBMid13), .HiOut(wRegInB13), .LoOut(wRegInA14) );
BubbleSort_Node #( 32 ) BSN2_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid14), .BIn(wBMid14), .HiOut(wRegInB14), .LoOut(wRegInA15) );
BubbleSort_Node #( 32 ) BSN2_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid15), .BIn(wBMid15), .HiOut(wRegInB15), .LoOut(wRegInA16) );
BubbleSort_Node #( 32 ) BSN2_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid16), .BIn(wBMid16), .HiOut(wRegInB16), .LoOut(wRegInA17) );
BubbleSort_Node #( 32 ) BSN2_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid17), .BIn(wBMid17), .HiOut(wRegInB17), .LoOut(wRegInA18) );
BubbleSort_Node #( 32 ) BSN2_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid18), .BIn(wBMid18), .HiOut(wRegInB18), .LoOut(wRegInA19) );
BubbleSort_Node #( 32 ) BSN2_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid19), .BIn(wBMid19), .HiOut(wRegInB19), .LoOut(wRegInA20) );
BubbleSort_Node #( 32 ) BSN2_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid20), .BIn(wBMid20), .HiOut(wRegInB20), .LoOut(wRegInA21) );
BubbleSort_Node #( 32 ) BSN2_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid21), .BIn(wBMid21), .HiOut(wRegInB21), .LoOut(wRegInA22) );
BubbleSort_Node #( 32 ) BSN2_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid22), .BIn(wBMid22), .HiOut(wRegInB22), .LoOut(wRegInA23) );
BubbleSort_Node #( 32 ) BSN2_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid23), .BIn(wBMid23), .HiOut(wRegInB23), .LoOut(wRegInA24) );
BubbleSort_Node #( 32 ) BSN2_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid24), .BIn(wBMid24), .HiOut(wRegInB24), .LoOut(wRegInA25) );
BubbleSort_Node #( 32 ) BSN2_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid25), .BIn(wBMid25), .HiOut(wRegInB25), .LoOut(wRegInA26) );
BubbleSort_Node #( 32 ) BSN2_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid26), .BIn(wBMid26), .HiOut(wRegInB26), .LoOut(wRegInA27) );
BubbleSort_Node #( 32 ) BSN2_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid27), .BIn(wBMid27), .HiOut(wRegInB27), .LoOut(wRegInA28) );
BubbleSort_Node #( 32 ) BSN2_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid28), .BIn(wBMid28), .HiOut(wRegInB28), .LoOut(wRegInA29) );
BubbleSort_Node #( 32 ) BSN2_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid29), .BIn(wBMid29), .HiOut(wRegInB29), .LoOut(wRegInA30) );
BubbleSort_Node #( 32 ) BSN2_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid30), .BIn(wBMid30), .HiOut(wRegInB30), .LoOut(wRegInA31) );
BubbleSort_Node #( 32 ) BSN2_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid31), .BIn(wBMid31), .HiOut(wRegInB31), .LoOut(wRegInA32) );
BubbleSort_Node #( 32 ) BSN2_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid32), .BIn(wBMid32), .HiOut(wRegInB32), .LoOut(wRegInA33) );
BubbleSort_Node #( 32 ) BSN2_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid33), .BIn(wBMid33), .HiOut(wRegInB33), .LoOut(wRegInA34) );
BubbleSort_Node #( 32 ) BSN2_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid34), .BIn(wBMid34), .HiOut(wRegInB34), .LoOut(wRegInA35) );
BubbleSort_Node #( 32 ) BSN2_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid35), .BIn(wBMid35), .HiOut(wRegInB35), .LoOut(wRegInA36) );
BubbleSort_Node #( 32 ) BSN2_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid36), .BIn(wBMid36), .HiOut(wRegInB36), .LoOut(wRegInA37) );
BubbleSort_Node #( 32 ) BSN2_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid37), .BIn(wBMid37), .HiOut(wRegInB37), .LoOut(wRegInA38) );
BubbleSort_Node #( 32 ) BSN2_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid38), .BIn(wBMid38), .HiOut(wRegInB38), .LoOut(wRegInA39) );
BubbleSort_Node #( 32 ) BSN2_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid39), .BIn(wBMid39), .HiOut(wRegInB39), .LoOut(wRegInA40) );
BubbleSort_Node #( 32 ) BSN2_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid40), .BIn(wBMid40), .HiOut(wRegInB40), .LoOut(wRegInA41) );
BubbleSort_Node #( 32 ) BSN2_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid41), .BIn(wBMid41), .HiOut(wRegInB41), .LoOut(wRegInA42) );
BubbleSort_Node #( 32 ) BSN2_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid42), .BIn(wBMid42), .HiOut(wRegInB42), .LoOut(wRegInA43) );
BubbleSort_Node #( 32 ) BSN2_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid43), .BIn(wBMid43), .HiOut(wRegInB43), .LoOut(wRegInA44) );
BubbleSort_Node #( 32 ) BSN2_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid44), .BIn(wBMid44), .HiOut(wRegInB44), .LoOut(wRegInA45) );
BubbleSort_Node #( 32 ) BSN2_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid45), .BIn(wBMid45), .HiOut(wRegInB45), .LoOut(wRegInA46) );
BubbleSort_Node #( 32 ) BSN2_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid46), .BIn(wBMid46), .HiOut(wRegInB46), .LoOut(wRegInA47) );
BubbleSort_Node #( 32 ) BSN2_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid47), .BIn(wBMid47), .HiOut(wRegInB47), .LoOut(wRegInA48) );
BubbleSort_Node #( 32 ) BSN2_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid48), .BIn(wBMid48), .HiOut(wRegInB48), .LoOut(wRegInA49) );
BubbleSort_Node #( 32 ) BSN2_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid49), .BIn(wBMid49), .HiOut(wRegInB49), .LoOut(wRegInA50) );
BubbleSort_Node #( 32 ) BSN2_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid50), .BIn(wBMid50), .HiOut(wRegInB50), .LoOut(wRegInA51) );
BubbleSort_Node #( 32 ) BSN2_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid51), .BIn(wBMid51), .HiOut(wRegInB51), .LoOut(wRegInA52) );
BubbleSort_Node #( 32 ) BSN2_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid52), .BIn(wBMid52), .HiOut(wRegInB52), .LoOut(wRegInA53) );
BubbleSort_Node #( 32 ) BSN2_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid53), .BIn(wBMid53), .HiOut(wRegInB53), .LoOut(wRegInA54) );
BubbleSort_Node #( 32 ) BSN2_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid54), .BIn(wBMid54), .HiOut(wRegInB54), .LoOut(wRegInA55) );
BubbleSort_Node #( 32 ) BSN2_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid55), .BIn(wBMid55), .HiOut(wRegInB55), .LoOut(wRegInA56) );
BubbleSort_Node #( 32 ) BSN2_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid56), .BIn(wBMid56), .HiOut(wRegInB56), .LoOut(wRegInA57) );
BubbleSort_Node #( 32 ) BSN2_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid57), .BIn(wBMid57), .HiOut(wRegInB57), .LoOut(wRegInA58) );
BubbleSort_Node #( 32 ) BSN2_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid58), .BIn(wBMid58), .HiOut(wRegInB58), .LoOut(wRegInA59) );
BubbleSort_Node #( 32 ) BSN2_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid59), .BIn(wBMid59), .HiOut(wRegInB59), .LoOut(wRegInA60) );
BubbleSort_Node #( 32 ) BSN2_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid60), .BIn(wBMid60), .HiOut(wRegInB60), .LoOut(wRegInA61) );
BubbleSort_Node #( 32 ) BSN2_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid61), .BIn(wBMid61), .HiOut(wRegInB61), .LoOut(wRegInA62) );
BubbleSort_Node #( 32 ) BSN2_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid62), .BIn(wBMid62), .HiOut(wRegInB62), .LoOut(wRegInA63) );
BubbleSort_Node #( 32 ) BSN2_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid63), .BIn(wBMid63), .HiOut(wRegInB63), .LoOut(wRegInA64) );
BubbleSort_Node #( 32 ) BSN2_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid64), .BIn(wBMid64), .HiOut(wRegInB64), .LoOut(wRegInA65) );
BubbleSort_Node #( 32 ) BSN2_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid65), .BIn(wBMid65), .HiOut(wRegInB65), .LoOut(wRegInA66) );
BubbleSort_Node #( 32 ) BSN2_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid66), .BIn(wBMid66), .HiOut(wRegInB66), .LoOut(wRegInA67) );
BubbleSort_Node #( 32 ) BSN2_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid67), .BIn(wBMid67), .HiOut(wRegInB67), .LoOut(wRegInA68) );
BubbleSort_Node #( 32 ) BSN2_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid68), .BIn(wBMid68), .HiOut(wRegInB68), .LoOut(wRegInA69) );
BubbleSort_Node #( 32 ) BSN2_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid69), .BIn(wBMid69), .HiOut(wRegInB69), .LoOut(wRegInA70) );
BubbleSort_Node #( 32 ) BSN2_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid70), .BIn(wBMid70), .HiOut(wRegInB70), .LoOut(wRegInA71) );
BubbleSort_Node #( 32 ) BSN2_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid71), .BIn(wBMid71), .HiOut(wRegInB71), .LoOut(wRegInA72) );
BubbleSort_Node #( 32 ) BSN2_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid72), .BIn(wBMid72), .HiOut(wRegInB72), .LoOut(wRegInA73) );
BubbleSort_Node #( 32 ) BSN2_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid73), .BIn(wBMid73), .HiOut(wRegInB73), .LoOut(wRegInA74) );
BubbleSort_Node #( 32 ) BSN2_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid74), .BIn(wBMid74), .HiOut(wRegInB74), .LoOut(wRegInA75) );
BubbleSort_Node #( 32 ) BSN2_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid75), .BIn(wBMid75), .HiOut(wRegInB75), .LoOut(wRegInA76) );
BubbleSort_Node #( 32 ) BSN2_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid76), .BIn(wBMid76), .HiOut(wRegInB76), .LoOut(wRegInA77) );
BubbleSort_Node #( 32 ) BSN2_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid77), .BIn(wBMid77), .HiOut(wRegInB77), .LoOut(wRegInA78) );
BubbleSort_Node #( 32 ) BSN2_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid78), .BIn(wBMid78), .HiOut(wRegInB78), .LoOut(wRegInA79) );
BubbleSort_Node #( 32 ) BSN2_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid79), .BIn(wBMid79), .HiOut(wRegInB79), .LoOut(wRegInA80) );
BubbleSort_Node #( 32 ) BSN2_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid80), .BIn(wBMid80), .HiOut(wRegInB80), .LoOut(wRegInA81) );
BubbleSort_Node #( 32 ) BSN2_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid81), .BIn(wBMid81), .HiOut(wRegInB81), .LoOut(wRegInA82) );
BubbleSort_Node #( 32 ) BSN2_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid82), .BIn(wBMid82), .HiOut(wRegInB82), .LoOut(wRegInA83) );
BubbleSort_Node #( 32 ) BSN2_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid83), .BIn(wBMid83), .HiOut(wRegInB83), .LoOut(wRegInA84) );
BubbleSort_Node #( 32 ) BSN2_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid84), .BIn(wBMid84), .HiOut(wRegInB84), .LoOut(wRegInA85) );
BubbleSort_Node #( 32 ) BSN2_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid85), .BIn(wBMid85), .HiOut(wRegInB85), .LoOut(wRegInA86) );
BubbleSort_Node #( 32 ) BSN2_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid86), .BIn(wBMid86), .HiOut(wRegInB86), .LoOut(wRegInA87) );
BubbleSort_Node #( 32 ) BSN2_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid87), .BIn(wBMid87), .HiOut(wRegInB87), .LoOut(wRegInA88) );
BubbleSort_Node #( 32 ) BSN2_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid88), .BIn(wBMid88), .HiOut(wRegInB88), .LoOut(wRegInA89) );
BubbleSort_Node #( 32 ) BSN2_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid89), .BIn(wBMid89), .HiOut(wRegInB89), .LoOut(wRegInA90) );
BubbleSort_Node #( 32 ) BSN2_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid90), .BIn(wBMid90), .HiOut(wRegInB90), .LoOut(wRegInA91) );
BubbleSort_Node #( 32 ) BSN2_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid91), .BIn(wBMid91), .HiOut(wRegInB91), .LoOut(wRegInA92) );
BubbleSort_Node #( 32 ) BSN2_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid92), .BIn(wBMid92), .HiOut(wRegInB92), .LoOut(wRegInA93) );
BubbleSort_Node #( 32 ) BSN2_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid93), .BIn(wBMid93), .HiOut(wRegInB93), .LoOut(wRegInA94) );
BubbleSort_Node #( 32 ) BSN2_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid94), .BIn(wBMid94), .HiOut(wRegInB94), .LoOut(wRegInA95) );
BubbleSort_Node #( 32 ) BSN2_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid95), .BIn(wBMid95), .HiOut(wRegInB95), .LoOut(wRegInA96) );
BubbleSort_Node #( 32 ) BSN2_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid96), .BIn(wBMid96), .HiOut(wRegInB96), .LoOut(wRegInA97) );
BubbleSort_Node #( 32 ) BSN2_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid97), .BIn(wBMid97), .HiOut(wRegInB97), .LoOut(wRegInA98) );
BubbleSort_Node #( 32 ) BSN2_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid98), .BIn(wBMid98), .HiOut(wRegInB98), .LoOut(wRegInA99) );
BubbleSort_Node #( 32 ) BSN2_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid99), .BIn(wBMid99), .HiOut(wRegInB99), .LoOut(wRegInA100) );
BubbleSort_Node #( 32 ) BSN2_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid100), .BIn(wBMid100), .HiOut(wRegInB100), .LoOut(wRegInA101) );
BubbleSort_Node #( 32 ) BSN2_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid101), .BIn(wBMid101), .HiOut(wRegInB101), .LoOut(wRegInA102) );
BubbleSort_Node #( 32 ) BSN2_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid102), .BIn(wBMid102), .HiOut(wRegInB102), .LoOut(wRegInA103) );
BubbleSort_Node #( 32 ) BSN2_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid103), .BIn(wBMid103), .HiOut(wRegInB103), .LoOut(wRegInA104) );
BubbleSort_Node #( 32 ) BSN2_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid104), .BIn(wBMid104), .HiOut(wRegInB104), .LoOut(wRegInA105) );
BubbleSort_Node #( 32 ) BSN2_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid105), .BIn(wBMid105), .HiOut(wRegInB105), .LoOut(wRegInA106) );
BubbleSort_Node #( 32 ) BSN2_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid106), .BIn(wBMid106), .HiOut(wRegInB106), .LoOut(wRegInA107) );
BubbleSort_Node #( 32 ) BSN2_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid107), .BIn(wBMid107), .HiOut(wRegInB107), .LoOut(wRegInA108) );
BubbleSort_Node #( 32 ) BSN2_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid108), .BIn(wBMid108), .HiOut(wRegInB108), .LoOut(wRegInA109) );
BubbleSort_Node #( 32 ) BSN2_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid109), .BIn(wBMid109), .HiOut(wRegInB109), .LoOut(wRegInA110) );
BubbleSort_Node #( 32 ) BSN2_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid110), .BIn(wBMid110), .HiOut(wRegInB110), .LoOut(wRegInA111) );
BubbleSort_Node #( 32 ) BSN2_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid111), .BIn(wBMid111), .HiOut(wRegInB111), .LoOut(wRegInA112) );
BubbleSort_Node #( 32 ) BSN2_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid112), .BIn(wBMid112), .HiOut(wRegInB112), .LoOut(wRegInA113) );
BubbleSort_Node #( 32 ) BSN2_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid113), .BIn(wBMid113), .HiOut(wRegInB113), .LoOut(wRegInA114) );
BubbleSort_Node #( 32 ) BSN2_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid114), .BIn(wBMid114), .HiOut(wRegInB114), .LoOut(wRegInA115) );
BubbleSort_Node #( 32 ) BSN2_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid115), .BIn(wBMid115), .HiOut(wRegInB115), .LoOut(wRegInA116) );
BubbleSort_Node #( 32 ) BSN2_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid116), .BIn(wBMid116), .HiOut(wRegInB116), .LoOut(wRegInA117) );
BubbleSort_Node #( 32 ) BSN2_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid117), .BIn(wBMid117), .HiOut(wRegInB117), .LoOut(wRegInA118) );
BubbleSort_Node #( 32 ) BSN2_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid118), .BIn(wBMid118), .HiOut(wRegInB118), .LoOut(wRegInA119) );
BubbleSort_Node #( 32 ) BSN2_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid119), .BIn(wBMid119), .HiOut(wRegInB119), .LoOut(wRegInA120) );
BubbleSort_Node #( 32 ) BSN2_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid120), .BIn(wBMid120), .HiOut(wRegInB120), .LoOut(wRegInA121) );
BubbleSort_Node #( 32 ) BSN2_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid121), .BIn(wBMid121), .HiOut(wRegInB121), .LoOut(wRegInA122) );
BubbleSort_Node #( 32 ) BSN2_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid122), .BIn(wBMid122), .HiOut(wRegInB122), .LoOut(wRegInA123) );
BubbleSort_Node #( 32 ) BSN2_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid123), .BIn(wBMid123), .HiOut(wRegInB123), .LoOut(wRegInA124) );
BubbleSort_Node #( 32 ) BSN2_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid124), .BIn(wBMid124), .HiOut(wRegInB124), .LoOut(wRegInA125) );
BubbleSort_Node #( 32 ) BSN2_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid125), .BIn(wBMid125), .HiOut(wRegInB125), .LoOut(wRegInA126) );
BubbleSort_Node #( 32 ) BSN2_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid126), .BIn(wBMid126), .HiOut(wRegInB126), .LoOut(wRegInA127) );
BubbleSort_Node #( 32 ) BSN2_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid127), .BIn(wBMid127), .HiOut(wRegInB127), .LoOut(wRegInA128) );
BubbleSort_Node #( 32 ) BSN2_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid128), .BIn(wBMid128), .HiOut(wRegInB128), .LoOut(wRegInA129) );
BubbleSort_Node #( 32 ) BSN2_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid129), .BIn(wBMid129), .HiOut(wRegInB129), .LoOut(wRegInA130) );
BubbleSort_Node #( 32 ) BSN2_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid130), .BIn(wBMid130), .HiOut(wRegInB130), .LoOut(wRegInA131) );
BubbleSort_Node #( 32 ) BSN2_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid131), .BIn(wBMid131), .HiOut(wRegInB131), .LoOut(wRegInA132) );
BubbleSort_Node #( 32 ) BSN2_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid132), .BIn(wBMid132), .HiOut(wRegInB132), .LoOut(wRegInA133) );
BubbleSort_Node #( 32 ) BSN2_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid133), .BIn(wBMid133), .HiOut(wRegInB133), .LoOut(wRegInA134) );
BubbleSort_Node #( 32 ) BSN2_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid134), .BIn(wBMid134), .HiOut(wRegInB134), .LoOut(wRegInA135) );
BubbleSort_Node #( 32 ) BSN2_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid135), .BIn(wBMid135), .HiOut(wRegInB135), .LoOut(wRegInA136) );
BubbleSort_Node #( 32 ) BSN2_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid136), .BIn(wBMid136), .HiOut(wRegInB136), .LoOut(wRegInA137) );
BubbleSort_Node #( 32 ) BSN2_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid137), .BIn(wBMid137), .HiOut(wRegInB137), .LoOut(wRegInA138) );
BubbleSort_Node #( 32 ) BSN2_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid138), .BIn(wBMid138), .HiOut(wRegInB138), .LoOut(wRegInA139) );
BubbleSort_Node #( 32 ) BSN2_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid139), .BIn(wBMid139), .HiOut(wRegInB139), .LoOut(wRegInA140) );
BubbleSort_Node #( 32 ) BSN2_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid140), .BIn(wBMid140), .HiOut(wRegInB140), .LoOut(wRegInA141) );
BubbleSort_Node #( 32 ) BSN2_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid141), .BIn(wBMid141), .HiOut(wRegInB141), .LoOut(wRegInA142) );
BubbleSort_Node #( 32 ) BSN2_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid142), .BIn(wBMid142), .HiOut(wRegInB142), .LoOut(wRegInA143) );
BubbleSort_Node #( 32 ) BSN2_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid143), .BIn(wBMid143), .HiOut(wRegInB143), .LoOut(wRegInA144) );
BubbleSort_Node #( 32 ) BSN2_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid144), .BIn(wBMid144), .HiOut(wRegInB144), .LoOut(wRegInA145) );
BubbleSort_Node #( 32 ) BSN2_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid145), .BIn(wBMid145), .HiOut(wRegInB145), .LoOut(wRegInA146) );
BubbleSort_Node #( 32 ) BSN2_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid146), .BIn(wBMid146), .HiOut(wRegInB146), .LoOut(wRegInA147) );
BubbleSort_Node #( 32 ) BSN2_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid147), .BIn(wBMid147), .HiOut(wRegInB147), .LoOut(wRegInA148) );
BubbleSort_Node #( 32 ) BSN2_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid148), .BIn(wBMid148), .HiOut(wRegInB148), .LoOut(wRegInA149) );
BubbleSort_Node #( 32 ) BSN2_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid149), .BIn(wBMid149), .HiOut(wRegInB149), .LoOut(wRegInA150) );
BubbleSort_Node #( 32 ) BSN2_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid150), .BIn(wBMid150), .HiOut(wRegInB150), .LoOut(wRegInA151) );
BubbleSort_Node #( 32 ) BSN2_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid151), .BIn(wBMid151), .HiOut(wRegInB151), .LoOut(wRegInA152) );
BubbleSort_Node #( 32 ) BSN2_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid152), .BIn(wBMid152), .HiOut(wRegInB152), .LoOut(wRegInA153) );
BubbleSort_Node #( 32 ) BSN2_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid153), .BIn(wBMid153), .HiOut(wRegInB153), .LoOut(wRegInA154) );
BubbleSort_Node #( 32 ) BSN2_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid154), .BIn(wBMid154), .HiOut(wRegInB154), .LoOut(wRegInA155) );
BubbleSort_Node #( 32 ) BSN2_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid155), .BIn(wBMid155), .HiOut(wRegInB155), .LoOut(wRegInA156) );
BubbleSort_Node #( 32 ) BSN2_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid156), .BIn(wBMid156), .HiOut(wRegInB156), .LoOut(wRegInA157) );
BubbleSort_Node #( 32 ) BSN2_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid157), .BIn(wBMid157), .HiOut(wRegInB157), .LoOut(wRegInA158) );
BubbleSort_Node #( 32 ) BSN2_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid158), .BIn(wBMid158), .HiOut(wRegInB158), .LoOut(wRegInA159) );
BubbleSort_Node #( 32 ) BSN2_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid159), .BIn(wBMid159), .HiOut(wRegInB159), .LoOut(wRegInA160) );
BubbleSort_Node #( 32 ) BSN2_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid160), .BIn(wBMid160), .HiOut(wRegInB160), .LoOut(wRegInA161) );
BubbleSort_Node #( 32 ) BSN2_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid161), .BIn(wBMid161), .HiOut(wRegInB161), .LoOut(wRegInA162) );
BubbleSort_Node #( 32 ) BSN2_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid162), .BIn(wBMid162), .HiOut(wRegInB162), .LoOut(wRegInA163) );
BubbleSort_Node #( 32 ) BSN2_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid163), .BIn(wBMid163), .HiOut(wRegInB163), .LoOut(wRegInA164) );
BubbleSort_Node #( 32 ) BSN2_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid164), .BIn(wBMid164), .HiOut(wRegInB164), .LoOut(wRegInA165) );
BubbleSort_Node #( 32 ) BSN2_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid165), .BIn(wBMid165), .HiOut(wRegInB165), .LoOut(wRegInA166) );
BubbleSort_Node #( 32 ) BSN2_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid166), .BIn(wBMid166), .HiOut(wRegInB166), .LoOut(wRegInA167) );
BubbleSort_Node #( 32 ) BSN2_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid167), .BIn(wBMid167), .HiOut(wRegInB167), .LoOut(wRegInA168) );
BubbleSort_Node #( 32 ) BSN2_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid168), .BIn(wBMid168), .HiOut(wRegInB168), .LoOut(wRegInA169) );
BubbleSort_Node #( 32 ) BSN2_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid169), .BIn(wBMid169), .HiOut(wRegInB169), .LoOut(wRegInA170) );
BubbleSort_Node #( 32 ) BSN2_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid170), .BIn(wBMid170), .HiOut(wRegInB170), .LoOut(wRegInA171) );
BubbleSort_Node #( 32 ) BSN2_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid171), .BIn(wBMid171), .HiOut(wRegInB171), .LoOut(wRegInA172) );
BubbleSort_Node #( 32 ) BSN2_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid172), .BIn(wBMid172), .HiOut(wRegInB172), .LoOut(wRegInA173) );
BubbleSort_Node #( 32 ) BSN2_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid173), .BIn(wBMid173), .HiOut(wRegInB173), .LoOut(wRegInA174) );
BubbleSort_Node #( 32 ) BSN2_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid174), .BIn(wBMid174), .HiOut(wRegInB174), .LoOut(wRegInA175) );
BubbleSort_Node #( 32 ) BSN2_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid175), .BIn(wBMid175), .HiOut(wRegInB175), .LoOut(wRegInA176) );
BubbleSort_Node #( 32 ) BSN2_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid176), .BIn(wBMid176), .HiOut(wRegInB176), .LoOut(wRegInA177) );
BubbleSort_Node #( 32 ) BSN2_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid177), .BIn(wBMid177), .HiOut(wRegInB177), .LoOut(wRegInA178) );
BubbleSort_Node #( 32 ) BSN2_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid178), .BIn(wBMid178), .HiOut(wRegInB178), .LoOut(wRegInA179) );
BubbleSort_Node #( 32 ) BSN2_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid179), .BIn(wBMid179), .HiOut(wRegInB179), .LoOut(wRegInA180) );
BubbleSort_Node #( 32 ) BSN2_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid180), .BIn(wBMid180), .HiOut(wRegInB180), .LoOut(wRegInA181) );
BubbleSort_Node #( 32 ) BSN2_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid181), .BIn(wBMid181), .HiOut(wRegInB181), .LoOut(wRegInA182) );
BubbleSort_Node #( 32 ) BSN2_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid182), .BIn(wBMid182), .HiOut(wRegInB182), .LoOut(wRegInA183) );
BubbleSort_Node #( 32 ) BSN2_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid183), .BIn(wBMid183), .HiOut(wRegInB183), .LoOut(wRegInA184) );
BubbleSort_Node #( 32 ) BSN2_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid184), .BIn(wBMid184), .HiOut(wRegInB184), .LoOut(wRegInA185) );
BubbleSort_Node #( 32 ) BSN2_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid185), .BIn(wBMid185), .HiOut(wRegInB185), .LoOut(wRegInA186) );
BubbleSort_Node #( 32 ) BSN2_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid186), .BIn(wBMid186), .HiOut(wRegInB186), .LoOut(wRegInA187) );
BubbleSort_Node #( 32 ) BSN2_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid187), .BIn(wBMid187), .HiOut(wRegInB187), .LoOut(wRegInA188) );
BubbleSort_Node #( 32 ) BSN2_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid188), .BIn(wBMid188), .HiOut(wRegInB188), .LoOut(wRegInA189) );
BubbleSort_Node #( 32 ) BSN2_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid189), .BIn(wBMid189), .HiOut(wRegInB189), .LoOut(wRegInA190) );
BubbleSort_Node #( 32 ) BSN2_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid190), .BIn(wBMid190), .HiOut(wRegInB190), .LoOut(wRegInA191) );
BubbleSort_Node #( 32 ) BSN2_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid191), .BIn(wBMid191), .HiOut(wRegInB191), .LoOut(wRegInA192) );
BubbleSort_Node #( 32 ) BSN2_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid192), .BIn(wBMid192), .HiOut(wRegInB192), .LoOut(wRegInA193) );
BubbleSort_Node #( 32 ) BSN2_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid193), .BIn(wBMid193), .HiOut(wRegInB193), .LoOut(wRegInA194) );
BubbleSort_Node #( 32 ) BSN2_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid194), .BIn(wBMid194), .HiOut(wRegInB194), .LoOut(wRegInA195) );
BubbleSort_Node #( 32 ) BSN2_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid195), .BIn(wBMid195), .HiOut(wRegInB195), .LoOut(wRegInA196) );
BubbleSort_Node #( 32 ) BSN2_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid196), .BIn(wBMid196), .HiOut(wRegInB196), .LoOut(wRegInA197) );
BubbleSort_Node #( 32 ) BSN2_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid197), .BIn(wBMid197), .HiOut(wRegInB197), .LoOut(wRegInA198) );
BubbleSort_Node #( 32 ) BSN2_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid198), .BIn(wBMid198), .HiOut(wRegInB198), .LoOut(wRegInA199) );
BubbleSort_Node #( 32 ) BSN2_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid199), .BIn(wBMid199), .HiOut(wRegInB199), .LoOut(wRegInA200) );
BubbleSort_Node #( 32 ) BSN2_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid200), .BIn(wBMid200), .HiOut(wRegInB200), .LoOut(wRegInA201) );
BubbleSort_Node #( 32 ) BSN2_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid201), .BIn(wBMid201), .HiOut(wRegInB201), .LoOut(wRegInA202) );
BubbleSort_Node #( 32 ) BSN2_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid202), .BIn(wBMid202), .HiOut(wRegInB202), .LoOut(wRegInA203) );
BubbleSort_Node #( 32 ) BSN2_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid203), .BIn(wBMid203), .HiOut(wRegInB203), .LoOut(wRegInA204) );
BubbleSort_Node #( 32 ) BSN2_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid204), .BIn(wBMid204), .HiOut(wRegInB204), .LoOut(wRegInA205) );
BubbleSort_Node #( 32 ) BSN2_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid205), .BIn(wBMid205), .HiOut(wRegInB205), .LoOut(wRegInA206) );
BubbleSort_Node #( 32 ) BSN2_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid206), .BIn(wBMid206), .HiOut(wRegInB206), .LoOut(wRegInA207) );
BubbleSort_Node #( 32 ) BSN2_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid207), .BIn(wBMid207), .HiOut(wRegInB207), .LoOut(wRegInA208) );
BubbleSort_Node #( 32 ) BSN2_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid208), .BIn(wBMid208), .HiOut(wRegInB208), .LoOut(wRegInA209) );
BubbleSort_Node #( 32 ) BSN2_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid209), .BIn(wBMid209), .HiOut(wRegInB209), .LoOut(wRegInA210) );
BubbleSort_Node #( 32 ) BSN2_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid210), .BIn(wBMid210), .HiOut(wRegInB210), .LoOut(wRegInA211) );
BubbleSort_Node #( 32 ) BSN2_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid211), .BIn(wBMid211), .HiOut(wRegInB211), .LoOut(wRegInA212) );
BubbleSort_Node #( 32 ) BSN2_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid212), .BIn(wBMid212), .HiOut(wRegInB212), .LoOut(wRegInA213) );
BubbleSort_Node #( 32 ) BSN2_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid213), .BIn(wBMid213), .HiOut(wRegInB213), .LoOut(wRegInA214) );
BubbleSort_Node #( 32 ) BSN2_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid214), .BIn(wBMid214), .HiOut(wRegInB214), .LoOut(wRegInA215) );
BubbleSort_Node #( 32 ) BSN2_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid215), .BIn(wBMid215), .HiOut(wRegInB215), .LoOut(wRegInA216) );
BubbleSort_Node #( 32 ) BSN2_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid216), .BIn(wBMid216), .HiOut(wRegInB216), .LoOut(wRegInA217) );
BubbleSort_Node #( 32 ) BSN2_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid217), .BIn(wBMid217), .HiOut(wRegInB217), .LoOut(wRegInA218) );
BubbleSort_Node #( 32 ) BSN2_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid218), .BIn(wBMid218), .HiOut(wRegInB218), .LoOut(wRegInA219) );
BubbleSort_Node #( 32 ) BSN2_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid219), .BIn(wBMid219), .HiOut(wRegInB219), .LoOut(wRegInA220) );
BubbleSort_Node #( 32 ) BSN2_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid220), .BIn(wBMid220), .HiOut(wRegInB220), .LoOut(wRegInA221) );
BubbleSort_Node #( 32 ) BSN2_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid221), .BIn(wBMid221), .HiOut(wRegInB221), .LoOut(wRegInA222) );
BubbleSort_Node #( 32 ) BSN2_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid222), .BIn(wBMid222), .HiOut(wRegInB222), .LoOut(wRegInA223) );
BubbleSort_Node #( 32 ) BSN2_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid223), .BIn(wBMid223), .HiOut(wRegInB223), .LoOut(wRegInA224) );
BubbleSort_Node #( 32 ) BSN2_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid224), .BIn(wBMid224), .HiOut(wRegInB224), .LoOut(wRegInA225) );
BubbleSort_Node #( 32 ) BSN2_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid225), .BIn(wBMid225), .HiOut(wRegInB225), .LoOut(wRegInA226) );
BubbleSort_Node #( 32 ) BSN2_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid226), .BIn(wBMid226), .HiOut(wRegInB226), .LoOut(wRegInA227) );
BubbleSort_Node #( 32 ) BSN2_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid227), .BIn(wBMid227), .HiOut(wRegInB227), .LoOut(wRegInA228) );
BubbleSort_Node #( 32 ) BSN2_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid228), .BIn(wBMid228), .HiOut(wRegInB228), .LoOut(wRegInA229) );
BubbleSort_Node #( 32 ) BSN2_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid229), .BIn(wBMid229), .HiOut(wRegInB229), .LoOut(wRegInA230) );
BubbleSort_Node #( 32 ) BSN2_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid230), .BIn(wBMid230), .HiOut(wRegInB230), .LoOut(wRegInA231) );
BubbleSort_Node #( 32 ) BSN2_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid231), .BIn(wBMid231), .HiOut(wRegInB231), .LoOut(wRegInA232) );
BubbleSort_Node #( 32 ) BSN2_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid232), .BIn(wBMid232), .HiOut(wRegInB232), .LoOut(wRegInA233) );
BubbleSort_Node #( 32 ) BSN2_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid233), .BIn(wBMid233), .HiOut(wRegInB233), .LoOut(wRegInA234) );
BubbleSort_Node #( 32 ) BSN2_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid234), .BIn(wBMid234), .HiOut(wRegInB234), .LoOut(wRegInA235) );
BubbleSort_Node #( 32 ) BSN2_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid235), .BIn(wBMid235), .HiOut(wRegInB235), .LoOut(wRegInA236) );
BubbleSort_Node #( 32 ) BSN2_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid236), .BIn(wBMid236), .HiOut(wRegInB236), .LoOut(wRegInA237) );
BubbleSort_Node #( 32 ) BSN2_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid237), .BIn(wBMid237), .HiOut(wRegInB237), .LoOut(wRegInA238) );
BubbleSort_Node #( 32 ) BSN2_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid238), .BIn(wBMid238), .HiOut(wRegInB238), .LoOut(wRegInA239) );
BubbleSort_Node #( 32 ) BSN2_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid239), .BIn(wBMid239), .HiOut(wRegInB239), .LoOut(wRegInA240) );
BubbleSort_Node #( 32 ) BSN2_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid240), .BIn(wBMid240), .HiOut(wRegInB240), .LoOut(wRegInA241) );
BubbleSort_Node #( 32 ) BSN2_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid241), .BIn(wBMid241), .HiOut(wRegInB241), .LoOut(wRegInA242) );
BubbleSort_Node #( 32 ) BSN2_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid242), .BIn(wBMid242), .HiOut(wRegInB242), .LoOut(wRegInA243) );
BubbleSort_Node #( 32 ) BSN2_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid243), .BIn(wBMid243), .HiOut(wRegInB243), .LoOut(wRegInA244) );
BubbleSort_Node #( 32 ) BSN2_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid244), .BIn(wBMid244), .HiOut(wRegInB244), .LoOut(wRegInA245) );
BubbleSort_Node #( 32 ) BSN2_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid245), .BIn(wBMid245), .HiOut(wRegInB245), .LoOut(wRegInA246) );
BubbleSort_Node #( 32 ) BSN2_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid246), .BIn(wBMid246), .HiOut(wRegInB246), .LoOut(wRegInA247) );
BubbleSort_Node #( 32 ) BSN2_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid247), .BIn(wBMid247), .HiOut(wRegInB247), .LoOut(wRegInA248) );
BubbleSort_Node #( 32 ) BSN2_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid248), .BIn(wBMid248), .HiOut(wRegInB248), .LoOut(wRegInA249) );
BubbleSort_Node #( 32 ) BSN2_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid249), .BIn(wBMid249), .HiOut(wRegInB249), .LoOut(wRegInA250) );
BubbleSort_Node #( 32 ) BSN2_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid250), .BIn(wBMid250), .HiOut(wRegInB250), .LoOut(wRegInA251) );
BubbleSort_Node #( 32 ) BSN2_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid251), .BIn(wBMid251), .HiOut(wRegInB251), .LoOut(wRegInA252) );
BubbleSort_Node #( 32 ) BSN2_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid252), .BIn(wBMid252), .HiOut(wRegInB252), .LoOut(wRegInA253) );
BubbleSort_Node #( 32 ) BSN2_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid253), .BIn(wBMid253), .HiOut(wRegInB253), .LoOut(wRegInA254) );
BubbleSort_Node #( 32 ) BSN2_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .AIn(wAMid254), .BIn(wBMid254), .HiOut(wRegInB254), .LoOut(wRegInA255) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_511 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA0), .Out(wAIn0), .ScanIn(ScanLink512), .ScanOut(ScanLink511), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_510 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB0), .Out(wBIn0), .ScanIn(ScanLink511), .ScanOut(ScanLink510), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_509 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA1), .Out(wAIn1), .ScanIn(ScanLink510), .ScanOut(ScanLink509), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_508 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB1), .Out(wBIn1), .ScanIn(ScanLink509), .ScanOut(ScanLink508), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_507 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA2), .Out(wAIn2), .ScanIn(ScanLink508), .ScanOut(ScanLink507), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_506 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB2), .Out(wBIn2), .ScanIn(ScanLink507), .ScanOut(ScanLink506), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_505 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA3), .Out(wAIn3), .ScanIn(ScanLink506), .ScanOut(ScanLink505), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_504 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB3), .Out(wBIn3), .ScanIn(ScanLink505), .ScanOut(ScanLink504), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_503 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA4), .Out(wAIn4), .ScanIn(ScanLink504), .ScanOut(ScanLink503), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_502 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB4), .Out(wBIn4), .ScanIn(ScanLink503), .ScanOut(ScanLink502), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_501 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA5), .Out(wAIn5), .ScanIn(ScanLink502), .ScanOut(ScanLink501), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_500 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB5), .Out(wBIn5), .ScanIn(ScanLink501), .ScanOut(ScanLink500), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_499 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA6), .Out(wAIn6), .ScanIn(ScanLink500), .ScanOut(ScanLink499), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_498 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB6), .Out(wBIn6), .ScanIn(ScanLink499), .ScanOut(ScanLink498), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_497 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA7), .Out(wAIn7), .ScanIn(ScanLink498), .ScanOut(ScanLink497), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_496 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB7), .Out(wBIn7), .ScanIn(ScanLink497), .ScanOut(ScanLink496), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_495 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA8), .Out(wAIn8), .ScanIn(ScanLink496), .ScanOut(ScanLink495), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_494 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB8), .Out(wBIn8), .ScanIn(ScanLink495), .ScanOut(ScanLink494), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_493 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA9), .Out(wAIn9), .ScanIn(ScanLink494), .ScanOut(ScanLink493), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_492 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB9), .Out(wBIn9), .ScanIn(ScanLink493), .ScanOut(ScanLink492), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_491 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA10), .Out(wAIn10), .ScanIn(ScanLink492), .ScanOut(ScanLink491), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_490 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB10), .Out(wBIn10), .ScanIn(ScanLink491), .ScanOut(ScanLink490), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_489 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA11), .Out(wAIn11), .ScanIn(ScanLink490), .ScanOut(ScanLink489), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_488 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB11), .Out(wBIn11), .ScanIn(ScanLink489), .ScanOut(ScanLink488), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_487 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA12), .Out(wAIn12), .ScanIn(ScanLink488), .ScanOut(ScanLink487), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_486 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB12), .Out(wBIn12), .ScanIn(ScanLink487), .ScanOut(ScanLink486), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_485 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA13), .Out(wAIn13), .ScanIn(ScanLink486), .ScanOut(ScanLink485), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_484 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB13), .Out(wBIn13), .ScanIn(ScanLink485), .ScanOut(ScanLink484), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_483 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA14), .Out(wAIn14), .ScanIn(ScanLink484), .ScanOut(ScanLink483), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_482 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB14), .Out(wBIn14), .ScanIn(ScanLink483), .ScanOut(ScanLink482), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_481 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA15), .Out(wAIn15), .ScanIn(ScanLink482), .ScanOut(ScanLink481), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_480 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB15), .Out(wBIn15), .ScanIn(ScanLink481), .ScanOut(ScanLink480), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_479 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA16), .Out(wAIn16), .ScanIn(ScanLink480), .ScanOut(ScanLink479), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_478 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB16), .Out(wBIn16), .ScanIn(ScanLink479), .ScanOut(ScanLink478), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_477 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA17), .Out(wAIn17), .ScanIn(ScanLink478), .ScanOut(ScanLink477), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_476 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB17), .Out(wBIn17), .ScanIn(ScanLink477), .ScanOut(ScanLink476), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_475 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA18), .Out(wAIn18), .ScanIn(ScanLink476), .ScanOut(ScanLink475), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_474 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB18), .Out(wBIn18), .ScanIn(ScanLink475), .ScanOut(ScanLink474), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_473 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA19), .Out(wAIn19), .ScanIn(ScanLink474), .ScanOut(ScanLink473), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_472 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB19), .Out(wBIn19), .ScanIn(ScanLink473), .ScanOut(ScanLink472), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_471 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA20), .Out(wAIn20), .ScanIn(ScanLink472), .ScanOut(ScanLink471), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_470 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB20), .Out(wBIn20), .ScanIn(ScanLink471), .ScanOut(ScanLink470), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_469 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA21), .Out(wAIn21), .ScanIn(ScanLink470), .ScanOut(ScanLink469), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_468 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB21), .Out(wBIn21), .ScanIn(ScanLink469), .ScanOut(ScanLink468), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_467 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA22), .Out(wAIn22), .ScanIn(ScanLink468), .ScanOut(ScanLink467), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_466 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB22), .Out(wBIn22), .ScanIn(ScanLink467), .ScanOut(ScanLink466), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_465 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA23), .Out(wAIn23), .ScanIn(ScanLink466), .ScanOut(ScanLink465), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_464 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB23), .Out(wBIn23), .ScanIn(ScanLink465), .ScanOut(ScanLink464), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_463 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA24), .Out(wAIn24), .ScanIn(ScanLink464), .ScanOut(ScanLink463), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_462 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB24), .Out(wBIn24), .ScanIn(ScanLink463), .ScanOut(ScanLink462), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_461 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA25), .Out(wAIn25), .ScanIn(ScanLink462), .ScanOut(ScanLink461), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_460 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB25), .Out(wBIn25), .ScanIn(ScanLink461), .ScanOut(ScanLink460), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_459 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA26), .Out(wAIn26), .ScanIn(ScanLink460), .ScanOut(ScanLink459), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_458 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB26), .Out(wBIn26), .ScanIn(ScanLink459), .ScanOut(ScanLink458), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_457 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA27), .Out(wAIn27), .ScanIn(ScanLink458), .ScanOut(ScanLink457), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_456 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB27), .Out(wBIn27), .ScanIn(ScanLink457), .ScanOut(ScanLink456), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_455 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA28), .Out(wAIn28), .ScanIn(ScanLink456), .ScanOut(ScanLink455), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_454 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB28), .Out(wBIn28), .ScanIn(ScanLink455), .ScanOut(ScanLink454), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_453 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA29), .Out(wAIn29), .ScanIn(ScanLink454), .ScanOut(ScanLink453), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_452 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB29), .Out(wBIn29), .ScanIn(ScanLink453), .ScanOut(ScanLink452), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_451 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA30), .Out(wAIn30), .ScanIn(ScanLink452), .ScanOut(ScanLink451), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_450 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB30), .Out(wBIn30), .ScanIn(ScanLink451), .ScanOut(ScanLink450), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_449 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA31), .Out(wAIn31), .ScanIn(ScanLink450), .ScanOut(ScanLink449), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_448 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB31), .Out(wBIn31), .ScanIn(ScanLink449), .ScanOut(ScanLink448), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_447 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA32), .Out(wAIn32), .ScanIn(ScanLink448), .ScanOut(ScanLink447), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_446 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB32), .Out(wBIn32), .ScanIn(ScanLink447), .ScanOut(ScanLink446), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_445 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA33), .Out(wAIn33), .ScanIn(ScanLink446), .ScanOut(ScanLink445), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_444 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB33), .Out(wBIn33), .ScanIn(ScanLink445), .ScanOut(ScanLink444), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_443 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA34), .Out(wAIn34), .ScanIn(ScanLink444), .ScanOut(ScanLink443), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_442 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB34), .Out(wBIn34), .ScanIn(ScanLink443), .ScanOut(ScanLink442), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_441 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA35), .Out(wAIn35), .ScanIn(ScanLink442), .ScanOut(ScanLink441), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_440 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB35), .Out(wBIn35), .ScanIn(ScanLink441), .ScanOut(ScanLink440), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_439 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA36), .Out(wAIn36), .ScanIn(ScanLink440), .ScanOut(ScanLink439), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_438 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB36), .Out(wBIn36), .ScanIn(ScanLink439), .ScanOut(ScanLink438), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_437 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA37), .Out(wAIn37), .ScanIn(ScanLink438), .ScanOut(ScanLink437), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_436 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB37), .Out(wBIn37), .ScanIn(ScanLink437), .ScanOut(ScanLink436), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_435 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA38), .Out(wAIn38), .ScanIn(ScanLink436), .ScanOut(ScanLink435), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_434 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB38), .Out(wBIn38), .ScanIn(ScanLink435), .ScanOut(ScanLink434), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_433 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA39), .Out(wAIn39), .ScanIn(ScanLink434), .ScanOut(ScanLink433), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_432 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB39), .Out(wBIn39), .ScanIn(ScanLink433), .ScanOut(ScanLink432), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_431 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA40), .Out(wAIn40), .ScanIn(ScanLink432), .ScanOut(ScanLink431), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_430 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB40), .Out(wBIn40), .ScanIn(ScanLink431), .ScanOut(ScanLink430), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_429 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA41), .Out(wAIn41), .ScanIn(ScanLink430), .ScanOut(ScanLink429), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_428 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB41), .Out(wBIn41), .ScanIn(ScanLink429), .ScanOut(ScanLink428), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_427 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA42), .Out(wAIn42), .ScanIn(ScanLink428), .ScanOut(ScanLink427), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_426 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB42), .Out(wBIn42), .ScanIn(ScanLink427), .ScanOut(ScanLink426), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_425 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA43), .Out(wAIn43), .ScanIn(ScanLink426), .ScanOut(ScanLink425), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_424 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB43), .Out(wBIn43), .ScanIn(ScanLink425), .ScanOut(ScanLink424), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_423 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA44), .Out(wAIn44), .ScanIn(ScanLink424), .ScanOut(ScanLink423), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_422 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB44), .Out(wBIn44), .ScanIn(ScanLink423), .ScanOut(ScanLink422), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_421 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA45), .Out(wAIn45), .ScanIn(ScanLink422), .ScanOut(ScanLink421), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_420 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB45), .Out(wBIn45), .ScanIn(ScanLink421), .ScanOut(ScanLink420), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_419 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA46), .Out(wAIn46), .ScanIn(ScanLink420), .ScanOut(ScanLink419), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_418 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB46), .Out(wBIn46), .ScanIn(ScanLink419), .ScanOut(ScanLink418), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_417 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA47), .Out(wAIn47), .ScanIn(ScanLink418), .ScanOut(ScanLink417), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_416 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB47), .Out(wBIn47), .ScanIn(ScanLink417), .ScanOut(ScanLink416), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_415 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA48), .Out(wAIn48), .ScanIn(ScanLink416), .ScanOut(ScanLink415), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_414 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB48), .Out(wBIn48), .ScanIn(ScanLink415), .ScanOut(ScanLink414), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_413 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA49), .Out(wAIn49), .ScanIn(ScanLink414), .ScanOut(ScanLink413), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_412 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB49), .Out(wBIn49), .ScanIn(ScanLink413), .ScanOut(ScanLink412), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_411 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA50), .Out(wAIn50), .ScanIn(ScanLink412), .ScanOut(ScanLink411), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_410 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB50), .Out(wBIn50), .ScanIn(ScanLink411), .ScanOut(ScanLink410), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_409 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA51), .Out(wAIn51), .ScanIn(ScanLink410), .ScanOut(ScanLink409), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_408 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB51), .Out(wBIn51), .ScanIn(ScanLink409), .ScanOut(ScanLink408), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_407 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA52), .Out(wAIn52), .ScanIn(ScanLink408), .ScanOut(ScanLink407), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_406 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB52), .Out(wBIn52), .ScanIn(ScanLink407), .ScanOut(ScanLink406), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_405 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA53), .Out(wAIn53), .ScanIn(ScanLink406), .ScanOut(ScanLink405), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_404 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB53), .Out(wBIn53), .ScanIn(ScanLink405), .ScanOut(ScanLink404), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_403 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA54), .Out(wAIn54), .ScanIn(ScanLink404), .ScanOut(ScanLink403), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_402 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB54), .Out(wBIn54), .ScanIn(ScanLink403), .ScanOut(ScanLink402), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_401 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA55), .Out(wAIn55), .ScanIn(ScanLink402), .ScanOut(ScanLink401), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_400 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB55), .Out(wBIn55), .ScanIn(ScanLink401), .ScanOut(ScanLink400), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_399 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA56), .Out(wAIn56), .ScanIn(ScanLink400), .ScanOut(ScanLink399), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_398 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB56), .Out(wBIn56), .ScanIn(ScanLink399), .ScanOut(ScanLink398), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_397 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA57), .Out(wAIn57), .ScanIn(ScanLink398), .ScanOut(ScanLink397), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_396 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB57), .Out(wBIn57), .ScanIn(ScanLink397), .ScanOut(ScanLink396), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_395 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA58), .Out(wAIn58), .ScanIn(ScanLink396), .ScanOut(ScanLink395), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_394 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB58), .Out(wBIn58), .ScanIn(ScanLink395), .ScanOut(ScanLink394), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_393 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA59), .Out(wAIn59), .ScanIn(ScanLink394), .ScanOut(ScanLink393), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_392 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB59), .Out(wBIn59), .ScanIn(ScanLink393), .ScanOut(ScanLink392), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_391 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA60), .Out(wAIn60), .ScanIn(ScanLink392), .ScanOut(ScanLink391), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_390 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB60), .Out(wBIn60), .ScanIn(ScanLink391), .ScanOut(ScanLink390), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_389 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA61), .Out(wAIn61), .ScanIn(ScanLink390), .ScanOut(ScanLink389), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_388 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB61), .Out(wBIn61), .ScanIn(ScanLink389), .ScanOut(ScanLink388), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_387 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA62), .Out(wAIn62), .ScanIn(ScanLink388), .ScanOut(ScanLink387), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_386 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB62), .Out(wBIn62), .ScanIn(ScanLink387), .ScanOut(ScanLink386), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_385 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA63), .Out(wAIn63), .ScanIn(ScanLink386), .ScanOut(ScanLink385), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_384 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB63), .Out(wBIn63), .ScanIn(ScanLink385), .ScanOut(ScanLink384), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_383 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA64), .Out(wAIn64), .ScanIn(ScanLink384), .ScanOut(ScanLink383), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_382 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB64), .Out(wBIn64), .ScanIn(ScanLink383), .ScanOut(ScanLink382), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_381 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA65), .Out(wAIn65), .ScanIn(ScanLink382), .ScanOut(ScanLink381), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_380 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB65), .Out(wBIn65), .ScanIn(ScanLink381), .ScanOut(ScanLink380), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_379 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA66), .Out(wAIn66), .ScanIn(ScanLink380), .ScanOut(ScanLink379), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_378 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB66), .Out(wBIn66), .ScanIn(ScanLink379), .ScanOut(ScanLink378), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_377 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA67), .Out(wAIn67), .ScanIn(ScanLink378), .ScanOut(ScanLink377), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_376 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB67), .Out(wBIn67), .ScanIn(ScanLink377), .ScanOut(ScanLink376), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_375 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA68), .Out(wAIn68), .ScanIn(ScanLink376), .ScanOut(ScanLink375), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_374 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB68), .Out(wBIn68), .ScanIn(ScanLink375), .ScanOut(ScanLink374), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_373 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA69), .Out(wAIn69), .ScanIn(ScanLink374), .ScanOut(ScanLink373), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_372 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB69), .Out(wBIn69), .ScanIn(ScanLink373), .ScanOut(ScanLink372), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_371 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA70), .Out(wAIn70), .ScanIn(ScanLink372), .ScanOut(ScanLink371), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_370 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB70), .Out(wBIn70), .ScanIn(ScanLink371), .ScanOut(ScanLink370), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_369 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA71), .Out(wAIn71), .ScanIn(ScanLink370), .ScanOut(ScanLink369), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_368 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB71), .Out(wBIn71), .ScanIn(ScanLink369), .ScanOut(ScanLink368), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_367 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA72), .Out(wAIn72), .ScanIn(ScanLink368), .ScanOut(ScanLink367), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_366 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB72), .Out(wBIn72), .ScanIn(ScanLink367), .ScanOut(ScanLink366), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_365 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA73), .Out(wAIn73), .ScanIn(ScanLink366), .ScanOut(ScanLink365), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_364 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB73), .Out(wBIn73), .ScanIn(ScanLink365), .ScanOut(ScanLink364), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_363 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA74), .Out(wAIn74), .ScanIn(ScanLink364), .ScanOut(ScanLink363), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_362 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB74), .Out(wBIn74), .ScanIn(ScanLink363), .ScanOut(ScanLink362), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_361 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA75), .Out(wAIn75), .ScanIn(ScanLink362), .ScanOut(ScanLink361), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_360 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB75), .Out(wBIn75), .ScanIn(ScanLink361), .ScanOut(ScanLink360), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_359 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA76), .Out(wAIn76), .ScanIn(ScanLink360), .ScanOut(ScanLink359), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_358 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB76), .Out(wBIn76), .ScanIn(ScanLink359), .ScanOut(ScanLink358), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_357 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA77), .Out(wAIn77), .ScanIn(ScanLink358), .ScanOut(ScanLink357), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_356 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB77), .Out(wBIn77), .ScanIn(ScanLink357), .ScanOut(ScanLink356), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_355 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA78), .Out(wAIn78), .ScanIn(ScanLink356), .ScanOut(ScanLink355), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_354 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB78), .Out(wBIn78), .ScanIn(ScanLink355), .ScanOut(ScanLink354), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_353 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA79), .Out(wAIn79), .ScanIn(ScanLink354), .ScanOut(ScanLink353), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_352 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB79), .Out(wBIn79), .ScanIn(ScanLink353), .ScanOut(ScanLink352), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_351 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA80), .Out(wAIn80), .ScanIn(ScanLink352), .ScanOut(ScanLink351), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_350 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB80), .Out(wBIn80), .ScanIn(ScanLink351), .ScanOut(ScanLink350), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_349 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA81), .Out(wAIn81), .ScanIn(ScanLink350), .ScanOut(ScanLink349), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_348 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB81), .Out(wBIn81), .ScanIn(ScanLink349), .ScanOut(ScanLink348), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_347 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA82), .Out(wAIn82), .ScanIn(ScanLink348), .ScanOut(ScanLink347), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_346 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB82), .Out(wBIn82), .ScanIn(ScanLink347), .ScanOut(ScanLink346), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_345 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA83), .Out(wAIn83), .ScanIn(ScanLink346), .ScanOut(ScanLink345), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_344 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB83), .Out(wBIn83), .ScanIn(ScanLink345), .ScanOut(ScanLink344), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_343 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA84), .Out(wAIn84), .ScanIn(ScanLink344), .ScanOut(ScanLink343), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_342 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB84), .Out(wBIn84), .ScanIn(ScanLink343), .ScanOut(ScanLink342), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_341 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA85), .Out(wAIn85), .ScanIn(ScanLink342), .ScanOut(ScanLink341), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_340 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB85), .Out(wBIn85), .ScanIn(ScanLink341), .ScanOut(ScanLink340), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_339 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA86), .Out(wAIn86), .ScanIn(ScanLink340), .ScanOut(ScanLink339), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_338 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB86), .Out(wBIn86), .ScanIn(ScanLink339), .ScanOut(ScanLink338), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_337 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA87), .Out(wAIn87), .ScanIn(ScanLink338), .ScanOut(ScanLink337), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_336 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB87), .Out(wBIn87), .ScanIn(ScanLink337), .ScanOut(ScanLink336), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_335 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA88), .Out(wAIn88), .ScanIn(ScanLink336), .ScanOut(ScanLink335), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_334 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB88), .Out(wBIn88), .ScanIn(ScanLink335), .ScanOut(ScanLink334), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_333 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA89), .Out(wAIn89), .ScanIn(ScanLink334), .ScanOut(ScanLink333), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_332 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB89), .Out(wBIn89), .ScanIn(ScanLink333), .ScanOut(ScanLink332), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_331 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA90), .Out(wAIn90), .ScanIn(ScanLink332), .ScanOut(ScanLink331), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_330 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB90), .Out(wBIn90), .ScanIn(ScanLink331), .ScanOut(ScanLink330), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_329 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA91), .Out(wAIn91), .ScanIn(ScanLink330), .ScanOut(ScanLink329), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_328 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB91), .Out(wBIn91), .ScanIn(ScanLink329), .ScanOut(ScanLink328), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_327 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA92), .Out(wAIn92), .ScanIn(ScanLink328), .ScanOut(ScanLink327), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_326 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB92), .Out(wBIn92), .ScanIn(ScanLink327), .ScanOut(ScanLink326), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_325 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA93), .Out(wAIn93), .ScanIn(ScanLink326), .ScanOut(ScanLink325), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_324 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB93), .Out(wBIn93), .ScanIn(ScanLink325), .ScanOut(ScanLink324), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_323 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA94), .Out(wAIn94), .ScanIn(ScanLink324), .ScanOut(ScanLink323), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_322 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB94), .Out(wBIn94), .ScanIn(ScanLink323), .ScanOut(ScanLink322), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_321 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA95), .Out(wAIn95), .ScanIn(ScanLink322), .ScanOut(ScanLink321), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_320 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB95), .Out(wBIn95), .ScanIn(ScanLink321), .ScanOut(ScanLink320), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_319 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA96), .Out(wAIn96), .ScanIn(ScanLink320), .ScanOut(ScanLink319), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_318 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB96), .Out(wBIn96), .ScanIn(ScanLink319), .ScanOut(ScanLink318), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_317 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA97), .Out(wAIn97), .ScanIn(ScanLink318), .ScanOut(ScanLink317), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_316 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB97), .Out(wBIn97), .ScanIn(ScanLink317), .ScanOut(ScanLink316), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_315 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA98), .Out(wAIn98), .ScanIn(ScanLink316), .ScanOut(ScanLink315), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_314 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB98), .Out(wBIn98), .ScanIn(ScanLink315), .ScanOut(ScanLink314), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_313 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA99), .Out(wAIn99), .ScanIn(ScanLink314), .ScanOut(ScanLink313), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_312 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB99), .Out(wBIn99), .ScanIn(ScanLink313), .ScanOut(ScanLink312), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_311 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA100), .Out(wAIn100), .ScanIn(ScanLink312), .ScanOut(ScanLink311), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_310 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB100), .Out(wBIn100), .ScanIn(ScanLink311), .ScanOut(ScanLink310), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_309 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA101), .Out(wAIn101), .ScanIn(ScanLink310), .ScanOut(ScanLink309), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_308 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB101), .Out(wBIn101), .ScanIn(ScanLink309), .ScanOut(ScanLink308), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_307 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA102), .Out(wAIn102), .ScanIn(ScanLink308), .ScanOut(ScanLink307), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_306 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB102), .Out(wBIn102), .ScanIn(ScanLink307), .ScanOut(ScanLink306), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_305 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA103), .Out(wAIn103), .ScanIn(ScanLink306), .ScanOut(ScanLink305), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_304 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB103), .Out(wBIn103), .ScanIn(ScanLink305), .ScanOut(ScanLink304), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_303 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA104), .Out(wAIn104), .ScanIn(ScanLink304), .ScanOut(ScanLink303), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_302 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB104), .Out(wBIn104), .ScanIn(ScanLink303), .ScanOut(ScanLink302), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_301 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA105), .Out(wAIn105), .ScanIn(ScanLink302), .ScanOut(ScanLink301), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_300 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB105), .Out(wBIn105), .ScanIn(ScanLink301), .ScanOut(ScanLink300), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_299 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA106), .Out(wAIn106), .ScanIn(ScanLink300), .ScanOut(ScanLink299), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_298 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB106), .Out(wBIn106), .ScanIn(ScanLink299), .ScanOut(ScanLink298), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_297 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA107), .Out(wAIn107), .ScanIn(ScanLink298), .ScanOut(ScanLink297), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_296 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB107), .Out(wBIn107), .ScanIn(ScanLink297), .ScanOut(ScanLink296), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_295 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA108), .Out(wAIn108), .ScanIn(ScanLink296), .ScanOut(ScanLink295), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_294 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB108), .Out(wBIn108), .ScanIn(ScanLink295), .ScanOut(ScanLink294), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_293 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA109), .Out(wAIn109), .ScanIn(ScanLink294), .ScanOut(ScanLink293), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_292 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB109), .Out(wBIn109), .ScanIn(ScanLink293), .ScanOut(ScanLink292), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_291 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA110), .Out(wAIn110), .ScanIn(ScanLink292), .ScanOut(ScanLink291), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_290 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB110), .Out(wBIn110), .ScanIn(ScanLink291), .ScanOut(ScanLink290), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_289 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA111), .Out(wAIn111), .ScanIn(ScanLink290), .ScanOut(ScanLink289), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_288 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB111), .Out(wBIn111), .ScanIn(ScanLink289), .ScanOut(ScanLink288), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_287 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA112), .Out(wAIn112), .ScanIn(ScanLink288), .ScanOut(ScanLink287), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_286 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB112), .Out(wBIn112), .ScanIn(ScanLink287), .ScanOut(ScanLink286), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_285 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA113), .Out(wAIn113), .ScanIn(ScanLink286), .ScanOut(ScanLink285), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_284 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB113), .Out(wBIn113), .ScanIn(ScanLink285), .ScanOut(ScanLink284), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_283 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA114), .Out(wAIn114), .ScanIn(ScanLink284), .ScanOut(ScanLink283), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_282 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB114), .Out(wBIn114), .ScanIn(ScanLink283), .ScanOut(ScanLink282), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_281 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA115), .Out(wAIn115), .ScanIn(ScanLink282), .ScanOut(ScanLink281), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_280 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB115), .Out(wBIn115), .ScanIn(ScanLink281), .ScanOut(ScanLink280), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_279 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA116), .Out(wAIn116), .ScanIn(ScanLink280), .ScanOut(ScanLink279), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_278 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB116), .Out(wBIn116), .ScanIn(ScanLink279), .ScanOut(ScanLink278), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_277 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA117), .Out(wAIn117), .ScanIn(ScanLink278), .ScanOut(ScanLink277), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_276 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB117), .Out(wBIn117), .ScanIn(ScanLink277), .ScanOut(ScanLink276), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_275 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA118), .Out(wAIn118), .ScanIn(ScanLink276), .ScanOut(ScanLink275), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_274 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB118), .Out(wBIn118), .ScanIn(ScanLink275), .ScanOut(ScanLink274), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_273 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA119), .Out(wAIn119), .ScanIn(ScanLink274), .ScanOut(ScanLink273), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_272 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB119), .Out(wBIn119), .ScanIn(ScanLink273), .ScanOut(ScanLink272), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_271 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA120), .Out(wAIn120), .ScanIn(ScanLink272), .ScanOut(ScanLink271), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_270 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB120), .Out(wBIn120), .ScanIn(ScanLink271), .ScanOut(ScanLink270), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_269 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA121), .Out(wAIn121), .ScanIn(ScanLink270), .ScanOut(ScanLink269), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_268 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB121), .Out(wBIn121), .ScanIn(ScanLink269), .ScanOut(ScanLink268), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_267 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA122), .Out(wAIn122), .ScanIn(ScanLink268), .ScanOut(ScanLink267), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_266 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB122), .Out(wBIn122), .ScanIn(ScanLink267), .ScanOut(ScanLink266), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_265 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA123), .Out(wAIn123), .ScanIn(ScanLink266), .ScanOut(ScanLink265), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_264 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB123), .Out(wBIn123), .ScanIn(ScanLink265), .ScanOut(ScanLink264), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_263 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA124), .Out(wAIn124), .ScanIn(ScanLink264), .ScanOut(ScanLink263), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_262 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB124), .Out(wBIn124), .ScanIn(ScanLink263), .ScanOut(ScanLink262), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_261 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA125), .Out(wAIn125), .ScanIn(ScanLink262), .ScanOut(ScanLink261), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_260 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB125), .Out(wBIn125), .ScanIn(ScanLink261), .ScanOut(ScanLink260), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_259 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA126), .Out(wAIn126), .ScanIn(ScanLink260), .ScanOut(ScanLink259), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_258 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB126), .Out(wBIn126), .ScanIn(ScanLink259), .ScanOut(ScanLink258), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_257 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA127), .Out(wAIn127), .ScanIn(ScanLink258), .ScanOut(ScanLink257), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_256 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB127), .Out(wBIn127), .ScanIn(ScanLink257), .ScanOut(ScanLink256), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA128), .Out(wAIn128), .ScanIn(ScanLink256), .ScanOut(ScanLink255), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB128), .Out(wBIn128), .ScanIn(ScanLink255), .ScanOut(ScanLink254), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA129), .Out(wAIn129), .ScanIn(ScanLink254), .ScanOut(ScanLink253), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB129), .Out(wBIn129), .ScanIn(ScanLink253), .ScanOut(ScanLink252), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA130), .Out(wAIn130), .ScanIn(ScanLink252), .ScanOut(ScanLink251), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB130), .Out(wBIn130), .ScanIn(ScanLink251), .ScanOut(ScanLink250), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA131), .Out(wAIn131), .ScanIn(ScanLink250), .ScanOut(ScanLink249), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB131), .Out(wBIn131), .ScanIn(ScanLink249), .ScanOut(ScanLink248), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA132), .Out(wAIn132), .ScanIn(ScanLink248), .ScanOut(ScanLink247), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB132), .Out(wBIn132), .ScanIn(ScanLink247), .ScanOut(ScanLink246), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA133), .Out(wAIn133), .ScanIn(ScanLink246), .ScanOut(ScanLink245), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB133), .Out(wBIn133), .ScanIn(ScanLink245), .ScanOut(ScanLink244), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA134), .Out(wAIn134), .ScanIn(ScanLink244), .ScanOut(ScanLink243), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB134), .Out(wBIn134), .ScanIn(ScanLink243), .ScanOut(ScanLink242), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA135), .Out(wAIn135), .ScanIn(ScanLink242), .ScanOut(ScanLink241), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB135), .Out(wBIn135), .ScanIn(ScanLink241), .ScanOut(ScanLink240), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA136), .Out(wAIn136), .ScanIn(ScanLink240), .ScanOut(ScanLink239), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB136), .Out(wBIn136), .ScanIn(ScanLink239), .ScanOut(ScanLink238), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA137), .Out(wAIn137), .ScanIn(ScanLink238), .ScanOut(ScanLink237), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB137), .Out(wBIn137), .ScanIn(ScanLink237), .ScanOut(ScanLink236), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA138), .Out(wAIn138), .ScanIn(ScanLink236), .ScanOut(ScanLink235), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB138), .Out(wBIn138), .ScanIn(ScanLink235), .ScanOut(ScanLink234), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA139), .Out(wAIn139), .ScanIn(ScanLink234), .ScanOut(ScanLink233), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB139), .Out(wBIn139), .ScanIn(ScanLink233), .ScanOut(ScanLink232), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA140), .Out(wAIn140), .ScanIn(ScanLink232), .ScanOut(ScanLink231), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB140), .Out(wBIn140), .ScanIn(ScanLink231), .ScanOut(ScanLink230), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA141), .Out(wAIn141), .ScanIn(ScanLink230), .ScanOut(ScanLink229), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB141), .Out(wBIn141), .ScanIn(ScanLink229), .ScanOut(ScanLink228), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA142), .Out(wAIn142), .ScanIn(ScanLink228), .ScanOut(ScanLink227), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB142), .Out(wBIn142), .ScanIn(ScanLink227), .ScanOut(ScanLink226), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA143), .Out(wAIn143), .ScanIn(ScanLink226), .ScanOut(ScanLink225), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB143), .Out(wBIn143), .ScanIn(ScanLink225), .ScanOut(ScanLink224), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA144), .Out(wAIn144), .ScanIn(ScanLink224), .ScanOut(ScanLink223), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB144), .Out(wBIn144), .ScanIn(ScanLink223), .ScanOut(ScanLink222), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA145), .Out(wAIn145), .ScanIn(ScanLink222), .ScanOut(ScanLink221), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB145), .Out(wBIn145), .ScanIn(ScanLink221), .ScanOut(ScanLink220), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA146), .Out(wAIn146), .ScanIn(ScanLink220), .ScanOut(ScanLink219), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB146), .Out(wBIn146), .ScanIn(ScanLink219), .ScanOut(ScanLink218), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA147), .Out(wAIn147), .ScanIn(ScanLink218), .ScanOut(ScanLink217), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB147), .Out(wBIn147), .ScanIn(ScanLink217), .ScanOut(ScanLink216), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA148), .Out(wAIn148), .ScanIn(ScanLink216), .ScanOut(ScanLink215), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB148), .Out(wBIn148), .ScanIn(ScanLink215), .ScanOut(ScanLink214), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA149), .Out(wAIn149), .ScanIn(ScanLink214), .ScanOut(ScanLink213), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB149), .Out(wBIn149), .ScanIn(ScanLink213), .ScanOut(ScanLink212), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA150), .Out(wAIn150), .ScanIn(ScanLink212), .ScanOut(ScanLink211), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB150), .Out(wBIn150), .ScanIn(ScanLink211), .ScanOut(ScanLink210), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA151), .Out(wAIn151), .ScanIn(ScanLink210), .ScanOut(ScanLink209), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB151), .Out(wBIn151), .ScanIn(ScanLink209), .ScanOut(ScanLink208), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA152), .Out(wAIn152), .ScanIn(ScanLink208), .ScanOut(ScanLink207), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB152), .Out(wBIn152), .ScanIn(ScanLink207), .ScanOut(ScanLink206), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA153), .Out(wAIn153), .ScanIn(ScanLink206), .ScanOut(ScanLink205), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB153), .Out(wBIn153), .ScanIn(ScanLink205), .ScanOut(ScanLink204), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA154), .Out(wAIn154), .ScanIn(ScanLink204), .ScanOut(ScanLink203), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB154), .Out(wBIn154), .ScanIn(ScanLink203), .ScanOut(ScanLink202), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA155), .Out(wAIn155), .ScanIn(ScanLink202), .ScanOut(ScanLink201), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB155), .Out(wBIn155), .ScanIn(ScanLink201), .ScanOut(ScanLink200), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA156), .Out(wAIn156), .ScanIn(ScanLink200), .ScanOut(ScanLink199), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB156), .Out(wBIn156), .ScanIn(ScanLink199), .ScanOut(ScanLink198), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA157), .Out(wAIn157), .ScanIn(ScanLink198), .ScanOut(ScanLink197), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB157), .Out(wBIn157), .ScanIn(ScanLink197), .ScanOut(ScanLink196), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA158), .Out(wAIn158), .ScanIn(ScanLink196), .ScanOut(ScanLink195), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB158), .Out(wBIn158), .ScanIn(ScanLink195), .ScanOut(ScanLink194), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA159), .Out(wAIn159), .ScanIn(ScanLink194), .ScanOut(ScanLink193), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB159), .Out(wBIn159), .ScanIn(ScanLink193), .ScanOut(ScanLink192), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA160), .Out(wAIn160), .ScanIn(ScanLink192), .ScanOut(ScanLink191), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB160), .Out(wBIn160), .ScanIn(ScanLink191), .ScanOut(ScanLink190), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA161), .Out(wAIn161), .ScanIn(ScanLink190), .ScanOut(ScanLink189), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB161), .Out(wBIn161), .ScanIn(ScanLink189), .ScanOut(ScanLink188), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA162), .Out(wAIn162), .ScanIn(ScanLink188), .ScanOut(ScanLink187), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB162), .Out(wBIn162), .ScanIn(ScanLink187), .ScanOut(ScanLink186), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA163), .Out(wAIn163), .ScanIn(ScanLink186), .ScanOut(ScanLink185), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB163), .Out(wBIn163), .ScanIn(ScanLink185), .ScanOut(ScanLink184), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA164), .Out(wAIn164), .ScanIn(ScanLink184), .ScanOut(ScanLink183), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB164), .Out(wBIn164), .ScanIn(ScanLink183), .ScanOut(ScanLink182), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA165), .Out(wAIn165), .ScanIn(ScanLink182), .ScanOut(ScanLink181), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB165), .Out(wBIn165), .ScanIn(ScanLink181), .ScanOut(ScanLink180), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA166), .Out(wAIn166), .ScanIn(ScanLink180), .ScanOut(ScanLink179), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB166), .Out(wBIn166), .ScanIn(ScanLink179), .ScanOut(ScanLink178), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA167), .Out(wAIn167), .ScanIn(ScanLink178), .ScanOut(ScanLink177), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB167), .Out(wBIn167), .ScanIn(ScanLink177), .ScanOut(ScanLink176), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA168), .Out(wAIn168), .ScanIn(ScanLink176), .ScanOut(ScanLink175), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB168), .Out(wBIn168), .ScanIn(ScanLink175), .ScanOut(ScanLink174), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA169), .Out(wAIn169), .ScanIn(ScanLink174), .ScanOut(ScanLink173), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB169), .Out(wBIn169), .ScanIn(ScanLink173), .ScanOut(ScanLink172), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA170), .Out(wAIn170), .ScanIn(ScanLink172), .ScanOut(ScanLink171), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB170), .Out(wBIn170), .ScanIn(ScanLink171), .ScanOut(ScanLink170), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA171), .Out(wAIn171), .ScanIn(ScanLink170), .ScanOut(ScanLink169), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB171), .Out(wBIn171), .ScanIn(ScanLink169), .ScanOut(ScanLink168), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA172), .Out(wAIn172), .ScanIn(ScanLink168), .ScanOut(ScanLink167), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB172), .Out(wBIn172), .ScanIn(ScanLink167), .ScanOut(ScanLink166), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA173), .Out(wAIn173), .ScanIn(ScanLink166), .ScanOut(ScanLink165), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB173), .Out(wBIn173), .ScanIn(ScanLink165), .ScanOut(ScanLink164), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA174), .Out(wAIn174), .ScanIn(ScanLink164), .ScanOut(ScanLink163), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB174), .Out(wBIn174), .ScanIn(ScanLink163), .ScanOut(ScanLink162), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA175), .Out(wAIn175), .ScanIn(ScanLink162), .ScanOut(ScanLink161), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB175), .Out(wBIn175), .ScanIn(ScanLink161), .ScanOut(ScanLink160), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA176), .Out(wAIn176), .ScanIn(ScanLink160), .ScanOut(ScanLink159), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB176), .Out(wBIn176), .ScanIn(ScanLink159), .ScanOut(ScanLink158), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA177), .Out(wAIn177), .ScanIn(ScanLink158), .ScanOut(ScanLink157), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB177), .Out(wBIn177), .ScanIn(ScanLink157), .ScanOut(ScanLink156), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA178), .Out(wAIn178), .ScanIn(ScanLink156), .ScanOut(ScanLink155), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB178), .Out(wBIn178), .ScanIn(ScanLink155), .ScanOut(ScanLink154), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA179), .Out(wAIn179), .ScanIn(ScanLink154), .ScanOut(ScanLink153), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB179), .Out(wBIn179), .ScanIn(ScanLink153), .ScanOut(ScanLink152), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA180), .Out(wAIn180), .ScanIn(ScanLink152), .ScanOut(ScanLink151), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB180), .Out(wBIn180), .ScanIn(ScanLink151), .ScanOut(ScanLink150), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA181), .Out(wAIn181), .ScanIn(ScanLink150), .ScanOut(ScanLink149), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB181), .Out(wBIn181), .ScanIn(ScanLink149), .ScanOut(ScanLink148), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA182), .Out(wAIn182), .ScanIn(ScanLink148), .ScanOut(ScanLink147), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB182), .Out(wBIn182), .ScanIn(ScanLink147), .ScanOut(ScanLink146), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA183), .Out(wAIn183), .ScanIn(ScanLink146), .ScanOut(ScanLink145), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB183), .Out(wBIn183), .ScanIn(ScanLink145), .ScanOut(ScanLink144), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA184), .Out(wAIn184), .ScanIn(ScanLink144), .ScanOut(ScanLink143), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB184), .Out(wBIn184), .ScanIn(ScanLink143), .ScanOut(ScanLink142), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA185), .Out(wAIn185), .ScanIn(ScanLink142), .ScanOut(ScanLink141), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB185), .Out(wBIn185), .ScanIn(ScanLink141), .ScanOut(ScanLink140), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA186), .Out(wAIn186), .ScanIn(ScanLink140), .ScanOut(ScanLink139), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB186), .Out(wBIn186), .ScanIn(ScanLink139), .ScanOut(ScanLink138), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA187), .Out(wAIn187), .ScanIn(ScanLink138), .ScanOut(ScanLink137), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB187), .Out(wBIn187), .ScanIn(ScanLink137), .ScanOut(ScanLink136), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA188), .Out(wAIn188), .ScanIn(ScanLink136), .ScanOut(ScanLink135), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB188), .Out(wBIn188), .ScanIn(ScanLink135), .ScanOut(ScanLink134), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA189), .Out(wAIn189), .ScanIn(ScanLink134), .ScanOut(ScanLink133), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB189), .Out(wBIn189), .ScanIn(ScanLink133), .ScanOut(ScanLink132), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA190), .Out(wAIn190), .ScanIn(ScanLink132), .ScanOut(ScanLink131), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB190), .Out(wBIn190), .ScanIn(ScanLink131), .ScanOut(ScanLink130), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA191), .Out(wAIn191), .ScanIn(ScanLink130), .ScanOut(ScanLink129), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB191), .Out(wBIn191), .ScanIn(ScanLink129), .ScanOut(ScanLink128), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA192), .Out(wAIn192), .ScanIn(ScanLink128), .ScanOut(ScanLink127), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB192), .Out(wBIn192), .ScanIn(ScanLink127), .ScanOut(ScanLink126), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA193), .Out(wAIn193), .ScanIn(ScanLink126), .ScanOut(ScanLink125), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB193), .Out(wBIn193), .ScanIn(ScanLink125), .ScanOut(ScanLink124), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA194), .Out(wAIn194), .ScanIn(ScanLink124), .ScanOut(ScanLink123), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB194), .Out(wBIn194), .ScanIn(ScanLink123), .ScanOut(ScanLink122), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA195), .Out(wAIn195), .ScanIn(ScanLink122), .ScanOut(ScanLink121), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB195), .Out(wBIn195), .ScanIn(ScanLink121), .ScanOut(ScanLink120), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA196), .Out(wAIn196), .ScanIn(ScanLink120), .ScanOut(ScanLink119), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB196), .Out(wBIn196), .ScanIn(ScanLink119), .ScanOut(ScanLink118), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA197), .Out(wAIn197), .ScanIn(ScanLink118), .ScanOut(ScanLink117), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB197), .Out(wBIn197), .ScanIn(ScanLink117), .ScanOut(ScanLink116), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA198), .Out(wAIn198), .ScanIn(ScanLink116), .ScanOut(ScanLink115), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB198), .Out(wBIn198), .ScanIn(ScanLink115), .ScanOut(ScanLink114), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA199), .Out(wAIn199), .ScanIn(ScanLink114), .ScanOut(ScanLink113), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB199), .Out(wBIn199), .ScanIn(ScanLink113), .ScanOut(ScanLink112), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA200), .Out(wAIn200), .ScanIn(ScanLink112), .ScanOut(ScanLink111), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB200), .Out(wBIn200), .ScanIn(ScanLink111), .ScanOut(ScanLink110), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA201), .Out(wAIn201), .ScanIn(ScanLink110), .ScanOut(ScanLink109), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB201), .Out(wBIn201), .ScanIn(ScanLink109), .ScanOut(ScanLink108), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA202), .Out(wAIn202), .ScanIn(ScanLink108), .ScanOut(ScanLink107), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB202), .Out(wBIn202), .ScanIn(ScanLink107), .ScanOut(ScanLink106), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA203), .Out(wAIn203), .ScanIn(ScanLink106), .ScanOut(ScanLink105), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB203), .Out(wBIn203), .ScanIn(ScanLink105), .ScanOut(ScanLink104), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA204), .Out(wAIn204), .ScanIn(ScanLink104), .ScanOut(ScanLink103), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB204), .Out(wBIn204), .ScanIn(ScanLink103), .ScanOut(ScanLink102), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA205), .Out(wAIn205), .ScanIn(ScanLink102), .ScanOut(ScanLink101), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB205), .Out(wBIn205), .ScanIn(ScanLink101), .ScanOut(ScanLink100), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA206), .Out(wAIn206), .ScanIn(ScanLink100), .ScanOut(ScanLink99), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB206), .Out(wBIn206), .ScanIn(ScanLink99), .ScanOut(ScanLink98), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA207), .Out(wAIn207), .ScanIn(ScanLink98), .ScanOut(ScanLink97), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB207), .Out(wBIn207), .ScanIn(ScanLink97), .ScanOut(ScanLink96), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA208), .Out(wAIn208), .ScanIn(ScanLink96), .ScanOut(ScanLink95), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB208), .Out(wBIn208), .ScanIn(ScanLink95), .ScanOut(ScanLink94), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA209), .Out(wAIn209), .ScanIn(ScanLink94), .ScanOut(ScanLink93), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB209), .Out(wBIn209), .ScanIn(ScanLink93), .ScanOut(ScanLink92), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA210), .Out(wAIn210), .ScanIn(ScanLink92), .ScanOut(ScanLink91), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB210), .Out(wBIn210), .ScanIn(ScanLink91), .ScanOut(ScanLink90), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA211), .Out(wAIn211), .ScanIn(ScanLink90), .ScanOut(ScanLink89), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB211), .Out(wBIn211), .ScanIn(ScanLink89), .ScanOut(ScanLink88), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA212), .Out(wAIn212), .ScanIn(ScanLink88), .ScanOut(ScanLink87), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB212), .Out(wBIn212), .ScanIn(ScanLink87), .ScanOut(ScanLink86), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA213), .Out(wAIn213), .ScanIn(ScanLink86), .ScanOut(ScanLink85), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB213), .Out(wBIn213), .ScanIn(ScanLink85), .ScanOut(ScanLink84), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA214), .Out(wAIn214), .ScanIn(ScanLink84), .ScanOut(ScanLink83), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB214), .Out(wBIn214), .ScanIn(ScanLink83), .ScanOut(ScanLink82), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA215), .Out(wAIn215), .ScanIn(ScanLink82), .ScanOut(ScanLink81), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB215), .Out(wBIn215), .ScanIn(ScanLink81), .ScanOut(ScanLink80), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA216), .Out(wAIn216), .ScanIn(ScanLink80), .ScanOut(ScanLink79), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB216), .Out(wBIn216), .ScanIn(ScanLink79), .ScanOut(ScanLink78), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA217), .Out(wAIn217), .ScanIn(ScanLink78), .ScanOut(ScanLink77), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB217), .Out(wBIn217), .ScanIn(ScanLink77), .ScanOut(ScanLink76), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA218), .Out(wAIn218), .ScanIn(ScanLink76), .ScanOut(ScanLink75), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB218), .Out(wBIn218), .ScanIn(ScanLink75), .ScanOut(ScanLink74), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA219), .Out(wAIn219), .ScanIn(ScanLink74), .ScanOut(ScanLink73), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB219), .Out(wBIn219), .ScanIn(ScanLink73), .ScanOut(ScanLink72), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA220), .Out(wAIn220), .ScanIn(ScanLink72), .ScanOut(ScanLink71), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB220), .Out(wBIn220), .ScanIn(ScanLink71), .ScanOut(ScanLink70), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA221), .Out(wAIn221), .ScanIn(ScanLink70), .ScanOut(ScanLink69), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB221), .Out(wBIn221), .ScanIn(ScanLink69), .ScanOut(ScanLink68), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA222), .Out(wAIn222), .ScanIn(ScanLink68), .ScanOut(ScanLink67), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB222), .Out(wBIn222), .ScanIn(ScanLink67), .ScanOut(ScanLink66), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA223), .Out(wAIn223), .ScanIn(ScanLink66), .ScanOut(ScanLink65), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB223), .Out(wBIn223), .ScanIn(ScanLink65), .ScanOut(ScanLink64), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA224), .Out(wAIn224), .ScanIn(ScanLink64), .ScanOut(ScanLink63), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB224), .Out(wBIn224), .ScanIn(ScanLink63), .ScanOut(ScanLink62), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA225), .Out(wAIn225), .ScanIn(ScanLink62), .ScanOut(ScanLink61), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB225), .Out(wBIn225), .ScanIn(ScanLink61), .ScanOut(ScanLink60), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA226), .Out(wAIn226), .ScanIn(ScanLink60), .ScanOut(ScanLink59), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB226), .Out(wBIn226), .ScanIn(ScanLink59), .ScanOut(ScanLink58), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA227), .Out(wAIn227), .ScanIn(ScanLink58), .ScanOut(ScanLink57), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB227), .Out(wBIn227), .ScanIn(ScanLink57), .ScanOut(ScanLink56), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA228), .Out(wAIn228), .ScanIn(ScanLink56), .ScanOut(ScanLink55), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB228), .Out(wBIn228), .ScanIn(ScanLink55), .ScanOut(ScanLink54), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA229), .Out(wAIn229), .ScanIn(ScanLink54), .ScanOut(ScanLink53), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB229), .Out(wBIn229), .ScanIn(ScanLink53), .ScanOut(ScanLink52), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA230), .Out(wAIn230), .ScanIn(ScanLink52), .ScanOut(ScanLink51), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB230), .Out(wBIn230), .ScanIn(ScanLink51), .ScanOut(ScanLink50), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA231), .Out(wAIn231), .ScanIn(ScanLink50), .ScanOut(ScanLink49), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB231), .Out(wBIn231), .ScanIn(ScanLink49), .ScanOut(ScanLink48), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA232), .Out(wAIn232), .ScanIn(ScanLink48), .ScanOut(ScanLink47), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB232), .Out(wBIn232), .ScanIn(ScanLink47), .ScanOut(ScanLink46), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA233), .Out(wAIn233), .ScanIn(ScanLink46), .ScanOut(ScanLink45), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB233), .Out(wBIn233), .ScanIn(ScanLink45), .ScanOut(ScanLink44), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA234), .Out(wAIn234), .ScanIn(ScanLink44), .ScanOut(ScanLink43), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB234), .Out(wBIn234), .ScanIn(ScanLink43), .ScanOut(ScanLink42), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA235), .Out(wAIn235), .ScanIn(ScanLink42), .ScanOut(ScanLink41), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB235), .Out(wBIn235), .ScanIn(ScanLink41), .ScanOut(ScanLink40), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA236), .Out(wAIn236), .ScanIn(ScanLink40), .ScanOut(ScanLink39), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB236), .Out(wBIn236), .ScanIn(ScanLink39), .ScanOut(ScanLink38), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA237), .Out(wAIn237), .ScanIn(ScanLink38), .ScanOut(ScanLink37), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB237), .Out(wBIn237), .ScanIn(ScanLink37), .ScanOut(ScanLink36), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA238), .Out(wAIn238), .ScanIn(ScanLink36), .ScanOut(ScanLink35), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB238), .Out(wBIn238), .ScanIn(ScanLink35), .ScanOut(ScanLink34), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA239), .Out(wAIn239), .ScanIn(ScanLink34), .ScanOut(ScanLink33), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB239), .Out(wBIn239), .ScanIn(ScanLink33), .ScanOut(ScanLink32), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA240), .Out(wAIn240), .ScanIn(ScanLink32), .ScanOut(ScanLink31), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB240), .Out(wBIn240), .ScanIn(ScanLink31), .ScanOut(ScanLink30), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA241), .Out(wAIn241), .ScanIn(ScanLink30), .ScanOut(ScanLink29), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB241), .Out(wBIn241), .ScanIn(ScanLink29), .ScanOut(ScanLink28), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA242), .Out(wAIn242), .ScanIn(ScanLink28), .ScanOut(ScanLink27), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB242), .Out(wBIn242), .ScanIn(ScanLink27), .ScanOut(ScanLink26), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA243), .Out(wAIn243), .ScanIn(ScanLink26), .ScanOut(ScanLink25), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB243), .Out(wBIn243), .ScanIn(ScanLink25), .ScanOut(ScanLink24), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA244), .Out(wAIn244), .ScanIn(ScanLink24), .ScanOut(ScanLink23), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB244), .Out(wBIn244), .ScanIn(ScanLink23), .ScanOut(ScanLink22), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA245), .Out(wAIn245), .ScanIn(ScanLink22), .ScanOut(ScanLink21), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB245), .Out(wBIn245), .ScanIn(ScanLink21), .ScanOut(ScanLink20), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA246), .Out(wAIn246), .ScanIn(ScanLink20), .ScanOut(ScanLink19), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB246), .Out(wBIn246), .ScanIn(ScanLink19), .ScanOut(ScanLink18), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA247), .Out(wAIn247), .ScanIn(ScanLink18), .ScanOut(ScanLink17), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB247), .Out(wBIn247), .ScanIn(ScanLink17), .ScanOut(ScanLink16), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA248), .Out(wAIn248), .ScanIn(ScanLink16), .ScanOut(ScanLink15), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB248), .Out(wBIn248), .ScanIn(ScanLink15), .ScanOut(ScanLink14), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA249), .Out(wAIn249), .ScanIn(ScanLink14), .ScanOut(ScanLink13), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB249), .Out(wBIn249), .ScanIn(ScanLink13), .ScanOut(ScanLink12), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA250), .Out(wAIn250), .ScanIn(ScanLink12), .ScanOut(ScanLink11), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB250), .Out(wBIn250), .ScanIn(ScanLink11), .ScanOut(ScanLink10), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA251), .Out(wAIn251), .ScanIn(ScanLink10), .ScanOut(ScanLink9), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB251), .Out(wBIn251), .ScanIn(ScanLink9), .ScanOut(ScanLink8), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA252), .Out(wAIn252), .ScanIn(ScanLink8), .ScanOut(ScanLink7), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB252), .Out(wBIn252), .ScanIn(ScanLink7), .ScanOut(ScanLink6), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA253), .Out(wAIn253), .ScanIn(ScanLink6), .ScanOut(ScanLink5), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB253), .Out(wBIn253), .ScanIn(ScanLink5), .ScanOut(ScanLink4), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA254), .Out(wAIn254), .ScanIn(ScanLink4), .ScanOut(ScanLink3), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB254), .Out(wBIn254), .ScanIn(ScanLink3), .ScanOut(ScanLink2), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInA255), .Out(wAIn255), .ScanIn(ScanLink2), .ScanOut(ScanLink1), .ScanEnable(ScanEnable) );
BubbleSort_Reg #( 32, 1, 1 ) U_BSR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(wEnable), .In(wRegInB255), .Out(wBIn255), .ScanIn(ScanLink1), .ScanOut(ScanLink0), .ScanEnable(ScanEnable) );
BubbleSort_Control #( 9, 1, 32, 1 ) U_BSC ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Enable(wEnable), .ScanIn(ScanLink0), .ScanOut(ScanLink512), .ScanEnable(ScanEnable), .ScanId(1'd0) );

/*
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
