

/*
 *
 * RAW Benchmark Suite main defines
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/bheap/src/library.v,v 1.4 1997/08/09 05:56:52 jbabb Exp $
 *
 * Library for Binary Heap Benchmark
 *
 * Authors: Elliot Waingold         (elliotw@lcs.mit.edu)
 *          Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 * BHeap_Node is the basic three-way compare node (fully combinational)
 */

module BHeap_Node(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		  Enable, P_WR, P_In, P_Out,
		  L_WR, L_In, L_Out, R_WR, R_In, R_Out);

   parameter			 WIDTH=8;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* local connections */

   input			 Enable;
   output			 P_WR;
   input [WIDTH-1:0]		 P_In;
   output [WIDTH-1:0]		 P_Out;
   output			 L_WR;
   input [WIDTH-1:0]		 L_In;
   output [WIDTH-1:0]		 L_Out;
   output			 R_WR;
   input [WIDTH-1:0]		 R_In;
   output [WIDTH-1:0]		 R_Out;

   assign L_WR = (Enable && (L_In > P_In) && (L_In >= R_In));
   assign R_WR = (Enable && (R_In > P_In) && (R_In > L_In));
   assign P_WR = (L_WR || R_WR);

   assign P_Out = L_WR ? L_In : (R_WR ? R_In : `GlobalDataHighZ);
   assign L_Out = L_WR ? P_In : `GlobalDataHighZ;
   assign R_Out = R_WR ? P_In : `GlobalDataHighZ;

endmodule

/*
 * BHeap_Reg is a register with two inputs and two enables
 */

module BHeap_Reg(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		 ScanIn, ScanOut, ScanEnable,
		 Id, Out, Enable1, Enable2, In1, In2);

   parameter			 WIDTH=8,
	     IDWIDTH=8,
	     SCAN=1;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;


   /* local connections */

   input [IDWIDTH-1:0]		 Id;
   output [WIDTH-1:0]		 Out;
   reg [WIDTH-1:0]		 Out;
   input			 Enable1;
   input			 Enable2;
   input [WIDTH-1:0]		 In1;
   input [WIDTH-1:0]		 In2;


   /* support reading of the node data value (non-scan only) */

   assign 	DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out : `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;

   always @(posedge Clk)
      begin


	 /* reset will initialize the entire array to zero */

	 if (Reset)
	    Out = 0;


	 /* support scan in */

	 else if  (SCAN && ScanEnable)
	    Out = ScanIn[WIDTH-1:0];


	 /* support writing of the node data value (non-scan only) */

	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0] == Id))
	    Out = DataIn[WIDTH-1:0];


	 /* heap operation */

	 else if (Enable1)
	    Out = In1;
	 else if (Enable2)
	    Out = In2;
      end
endmodule


/*
 * BHeap_CtrlReg is a one-bit register used in shifting control from
 * level to level
 */

module BHeap_CtrlReg(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		     In, Out, Enable);

   parameter			 WIDTH=8;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* local connections */

   input			 In;
   output			 Out;
   reg				 Out;
   output			 Enable;

   assign Enable = Out;

   always @(posedge Clk)
      begin
	 if (Reset)
	    Out = 0;
	 else
	    Out = In;
      end
endmodule


/*
 * BHeap_Control is the controller node
 */

module BHeap_Control(Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		     ScanIn, ScanOut, ScanEnable, ScanId,
		     Id, Go, Done);

   parameter			 CWIDTH=8,
				 IDWIDTH=8,
				 WIDTH=8,
				 SCAN=1;


   /* global connections */

   input			 Clk, Reset, RD, WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;
   input [IDWIDTH-1:0]		 ScanId;


   /* local connections */

   input [IDWIDTH-1:0]		 Id;
   output			 Go;
   reg				 Go;
   input			 Done;


   /* a register for the counter and scan */

   reg [CWIDTH-1:0]		 Count;
   reg [WIDTH-1:0]		 ScanReg;


   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? Count :
         (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;

   always @(posedge Clk)
      begin
	 ScanReg = ScanIn;

	 Go = 0;
	 if (Reset)
	    begin
	       Count = 0;
	    end
	 else if (WR && (Addr[IDWIDTH-1:0] == Id))
	    begin
	       Count = DataIn[CWIDTH-1:0];
	       if (Count)
		  Go = 1;
	    end
	 else if (Done)
	    begin
	       Count = Count-1;
	       if (Count)
		  Go = 1;
	    end
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [0:0] wCtrlOut_0;
wire [0:0] wEnable_0;
wire [31:0] wRegInBot_0_0;
wire [0:0] wRegEnBot_0_0;
wire [31:0] wRegOut_0_0;
wire [0:0] wCtrlOut_1;
wire [0:0] wEnable_1;
wire [31:0] wRegInTop_1_0;
wire [0:0] wRegEnTop_1_0;
wire [31:0] wRegInBot_1_0;
wire [0:0] wRegEnBot_1_0;
wire [31:0] wRegOut_1_0;
wire [31:0] wRegInTop_1_1;
wire [0:0] wRegEnTop_1_1;
wire [31:0] wRegInBot_1_1;
wire [0:0] wRegEnBot_1_1;
wire [31:0] wRegOut_1_1;
wire [0:0] wCtrlOut_2;
wire [0:0] wEnable_2;
wire [31:0] wRegInTop_2_0;
wire [0:0] wRegEnTop_2_0;
wire [31:0] wRegInBot_2_0;
wire [0:0] wRegEnBot_2_0;
wire [31:0] wRegOut_2_0;
wire [31:0] wRegInTop_2_1;
wire [0:0] wRegEnTop_2_1;
wire [31:0] wRegInBot_2_1;
wire [0:0] wRegEnBot_2_1;
wire [31:0] wRegOut_2_1;
wire [31:0] wRegInTop_2_2;
wire [0:0] wRegEnTop_2_2;
wire [31:0] wRegInBot_2_2;
wire [0:0] wRegEnBot_2_2;
wire [31:0] wRegOut_2_2;
wire [31:0] wRegInTop_2_3;
wire [0:0] wRegEnTop_2_3;
wire [31:0] wRegInBot_2_3;
wire [0:0] wRegEnBot_2_3;
wire [31:0] wRegOut_2_3;
wire [0:0] wCtrlOut_3;
wire [0:0] wEnable_3;
wire [31:0] wRegInTop_3_0;
wire [0:0] wRegEnTop_3_0;
wire [31:0] wRegInBot_3_0;
wire [0:0] wRegEnBot_3_0;
wire [31:0] wRegOut_3_0;
wire [31:0] wRegInTop_3_1;
wire [0:0] wRegEnTop_3_1;
wire [31:0] wRegInBot_3_1;
wire [0:0] wRegEnBot_3_1;
wire [31:0] wRegOut_3_1;
wire [31:0] wRegInTop_3_2;
wire [0:0] wRegEnTop_3_2;
wire [31:0] wRegInBot_3_2;
wire [0:0] wRegEnBot_3_2;
wire [31:0] wRegOut_3_2;
wire [31:0] wRegInTop_3_3;
wire [0:0] wRegEnTop_3_3;
wire [31:0] wRegInBot_3_3;
wire [0:0] wRegEnBot_3_3;
wire [31:0] wRegOut_3_3;
wire [31:0] wRegInTop_3_4;
wire [0:0] wRegEnTop_3_4;
wire [31:0] wRegInBot_3_4;
wire [0:0] wRegEnBot_3_4;
wire [31:0] wRegOut_3_4;
wire [31:0] wRegInTop_3_5;
wire [0:0] wRegEnTop_3_5;
wire [31:0] wRegInBot_3_5;
wire [0:0] wRegEnBot_3_5;
wire [31:0] wRegOut_3_5;
wire [31:0] wRegInTop_3_6;
wire [0:0] wRegEnTop_3_6;
wire [31:0] wRegInBot_3_6;
wire [0:0] wRegEnBot_3_6;
wire [31:0] wRegOut_3_6;
wire [31:0] wRegInTop_3_7;
wire [0:0] wRegEnTop_3_7;
wire [31:0] wRegInBot_3_7;
wire [0:0] wRegEnBot_3_7;
wire [31:0] wRegOut_3_7;
wire [0:0] wCtrlOut_4;
wire [0:0] wEnable_4;
wire [31:0] wRegInTop_4_0;
wire [0:0] wRegEnTop_4_0;
wire [31:0] wRegInBot_4_0;
wire [0:0] wRegEnBot_4_0;
wire [31:0] wRegOut_4_0;
wire [31:0] wRegInTop_4_1;
wire [0:0] wRegEnTop_4_1;
wire [31:0] wRegInBot_4_1;
wire [0:0] wRegEnBot_4_1;
wire [31:0] wRegOut_4_1;
wire [31:0] wRegInTop_4_2;
wire [0:0] wRegEnTop_4_2;
wire [31:0] wRegInBot_4_2;
wire [0:0] wRegEnBot_4_2;
wire [31:0] wRegOut_4_2;
wire [31:0] wRegInTop_4_3;
wire [0:0] wRegEnTop_4_3;
wire [31:0] wRegInBot_4_3;
wire [0:0] wRegEnBot_4_3;
wire [31:0] wRegOut_4_3;
wire [31:0] wRegInTop_4_4;
wire [0:0] wRegEnTop_4_4;
wire [31:0] wRegInBot_4_4;
wire [0:0] wRegEnBot_4_4;
wire [31:0] wRegOut_4_4;
wire [31:0] wRegInTop_4_5;
wire [0:0] wRegEnTop_4_5;
wire [31:0] wRegInBot_4_5;
wire [0:0] wRegEnBot_4_5;
wire [31:0] wRegOut_4_5;
wire [31:0] wRegInTop_4_6;
wire [0:0] wRegEnTop_4_6;
wire [31:0] wRegInBot_4_6;
wire [0:0] wRegEnBot_4_6;
wire [31:0] wRegOut_4_6;
wire [31:0] wRegInTop_4_7;
wire [0:0] wRegEnTop_4_7;
wire [31:0] wRegInBot_4_7;
wire [0:0] wRegEnBot_4_7;
wire [31:0] wRegOut_4_7;
wire [31:0] wRegInTop_4_8;
wire [0:0] wRegEnTop_4_8;
wire [31:0] wRegInBot_4_8;
wire [0:0] wRegEnBot_4_8;
wire [31:0] wRegOut_4_8;
wire [31:0] wRegInTop_4_9;
wire [0:0] wRegEnTop_4_9;
wire [31:0] wRegInBot_4_9;
wire [0:0] wRegEnBot_4_9;
wire [31:0] wRegOut_4_9;
wire [31:0] wRegInTop_4_10;
wire [0:0] wRegEnTop_4_10;
wire [31:0] wRegInBot_4_10;
wire [0:0] wRegEnBot_4_10;
wire [31:0] wRegOut_4_10;
wire [31:0] wRegInTop_4_11;
wire [0:0] wRegEnTop_4_11;
wire [31:0] wRegInBot_4_11;
wire [0:0] wRegEnBot_4_11;
wire [31:0] wRegOut_4_11;
wire [31:0] wRegInTop_4_12;
wire [0:0] wRegEnTop_4_12;
wire [31:0] wRegInBot_4_12;
wire [0:0] wRegEnBot_4_12;
wire [31:0] wRegOut_4_12;
wire [31:0] wRegInTop_4_13;
wire [0:0] wRegEnTop_4_13;
wire [31:0] wRegInBot_4_13;
wire [0:0] wRegEnBot_4_13;
wire [31:0] wRegOut_4_13;
wire [31:0] wRegInTop_4_14;
wire [0:0] wRegEnTop_4_14;
wire [31:0] wRegInBot_4_14;
wire [0:0] wRegEnBot_4_14;
wire [31:0] wRegOut_4_14;
wire [31:0] wRegInTop_4_15;
wire [0:0] wRegEnTop_4_15;
wire [31:0] wRegInBot_4_15;
wire [0:0] wRegEnBot_4_15;
wire [31:0] wRegOut_4_15;
wire [0:0] wCtrlOut_5;
wire [0:0] wEnable_5;
wire [31:0] wRegInTop_5_0;
wire [0:0] wRegEnTop_5_0;
wire [31:0] wRegInBot_5_0;
wire [0:0] wRegEnBot_5_0;
wire [31:0] wRegOut_5_0;
wire [31:0] wRegInTop_5_1;
wire [0:0] wRegEnTop_5_1;
wire [31:0] wRegInBot_5_1;
wire [0:0] wRegEnBot_5_1;
wire [31:0] wRegOut_5_1;
wire [31:0] wRegInTop_5_2;
wire [0:0] wRegEnTop_5_2;
wire [31:0] wRegInBot_5_2;
wire [0:0] wRegEnBot_5_2;
wire [31:0] wRegOut_5_2;
wire [31:0] wRegInTop_5_3;
wire [0:0] wRegEnTop_5_3;
wire [31:0] wRegInBot_5_3;
wire [0:0] wRegEnBot_5_3;
wire [31:0] wRegOut_5_3;
wire [31:0] wRegInTop_5_4;
wire [0:0] wRegEnTop_5_4;
wire [31:0] wRegInBot_5_4;
wire [0:0] wRegEnBot_5_4;
wire [31:0] wRegOut_5_4;
wire [31:0] wRegInTop_5_5;
wire [0:0] wRegEnTop_5_5;
wire [31:0] wRegInBot_5_5;
wire [0:0] wRegEnBot_5_5;
wire [31:0] wRegOut_5_5;
wire [31:0] wRegInTop_5_6;
wire [0:0] wRegEnTop_5_6;
wire [31:0] wRegInBot_5_6;
wire [0:0] wRegEnBot_5_6;
wire [31:0] wRegOut_5_6;
wire [31:0] wRegInTop_5_7;
wire [0:0] wRegEnTop_5_7;
wire [31:0] wRegInBot_5_7;
wire [0:0] wRegEnBot_5_7;
wire [31:0] wRegOut_5_7;
wire [31:0] wRegInTop_5_8;
wire [0:0] wRegEnTop_5_8;
wire [31:0] wRegInBot_5_8;
wire [0:0] wRegEnBot_5_8;
wire [31:0] wRegOut_5_8;
wire [31:0] wRegInTop_5_9;
wire [0:0] wRegEnTop_5_9;
wire [31:0] wRegInBot_5_9;
wire [0:0] wRegEnBot_5_9;
wire [31:0] wRegOut_5_9;
wire [31:0] wRegInTop_5_10;
wire [0:0] wRegEnTop_5_10;
wire [31:0] wRegInBot_5_10;
wire [0:0] wRegEnBot_5_10;
wire [31:0] wRegOut_5_10;
wire [31:0] wRegInTop_5_11;
wire [0:0] wRegEnTop_5_11;
wire [31:0] wRegInBot_5_11;
wire [0:0] wRegEnBot_5_11;
wire [31:0] wRegOut_5_11;
wire [31:0] wRegInTop_5_12;
wire [0:0] wRegEnTop_5_12;
wire [31:0] wRegInBot_5_12;
wire [0:0] wRegEnBot_5_12;
wire [31:0] wRegOut_5_12;
wire [31:0] wRegInTop_5_13;
wire [0:0] wRegEnTop_5_13;
wire [31:0] wRegInBot_5_13;
wire [0:0] wRegEnBot_5_13;
wire [31:0] wRegOut_5_13;
wire [31:0] wRegInTop_5_14;
wire [0:0] wRegEnTop_5_14;
wire [31:0] wRegInBot_5_14;
wire [0:0] wRegEnBot_5_14;
wire [31:0] wRegOut_5_14;
wire [31:0] wRegInTop_5_15;
wire [0:0] wRegEnTop_5_15;
wire [31:0] wRegInBot_5_15;
wire [0:0] wRegEnBot_5_15;
wire [31:0] wRegOut_5_15;
wire [31:0] wRegInTop_5_16;
wire [0:0] wRegEnTop_5_16;
wire [31:0] wRegInBot_5_16;
wire [0:0] wRegEnBot_5_16;
wire [31:0] wRegOut_5_16;
wire [31:0] wRegInTop_5_17;
wire [0:0] wRegEnTop_5_17;
wire [31:0] wRegInBot_5_17;
wire [0:0] wRegEnBot_5_17;
wire [31:0] wRegOut_5_17;
wire [31:0] wRegInTop_5_18;
wire [0:0] wRegEnTop_5_18;
wire [31:0] wRegInBot_5_18;
wire [0:0] wRegEnBot_5_18;
wire [31:0] wRegOut_5_18;
wire [31:0] wRegInTop_5_19;
wire [0:0] wRegEnTop_5_19;
wire [31:0] wRegInBot_5_19;
wire [0:0] wRegEnBot_5_19;
wire [31:0] wRegOut_5_19;
wire [31:0] wRegInTop_5_20;
wire [0:0] wRegEnTop_5_20;
wire [31:0] wRegInBot_5_20;
wire [0:0] wRegEnBot_5_20;
wire [31:0] wRegOut_5_20;
wire [31:0] wRegInTop_5_21;
wire [0:0] wRegEnTop_5_21;
wire [31:0] wRegInBot_5_21;
wire [0:0] wRegEnBot_5_21;
wire [31:0] wRegOut_5_21;
wire [31:0] wRegInTop_5_22;
wire [0:0] wRegEnTop_5_22;
wire [31:0] wRegInBot_5_22;
wire [0:0] wRegEnBot_5_22;
wire [31:0] wRegOut_5_22;
wire [31:0] wRegInTop_5_23;
wire [0:0] wRegEnTop_5_23;
wire [31:0] wRegInBot_5_23;
wire [0:0] wRegEnBot_5_23;
wire [31:0] wRegOut_5_23;
wire [31:0] wRegInTop_5_24;
wire [0:0] wRegEnTop_5_24;
wire [31:0] wRegInBot_5_24;
wire [0:0] wRegEnBot_5_24;
wire [31:0] wRegOut_5_24;
wire [31:0] wRegInTop_5_25;
wire [0:0] wRegEnTop_5_25;
wire [31:0] wRegInBot_5_25;
wire [0:0] wRegEnBot_5_25;
wire [31:0] wRegOut_5_25;
wire [31:0] wRegInTop_5_26;
wire [0:0] wRegEnTop_5_26;
wire [31:0] wRegInBot_5_26;
wire [0:0] wRegEnBot_5_26;
wire [31:0] wRegOut_5_26;
wire [31:0] wRegInTop_5_27;
wire [0:0] wRegEnTop_5_27;
wire [31:0] wRegInBot_5_27;
wire [0:0] wRegEnBot_5_27;
wire [31:0] wRegOut_5_27;
wire [31:0] wRegInTop_5_28;
wire [0:0] wRegEnTop_5_28;
wire [31:0] wRegInBot_5_28;
wire [0:0] wRegEnBot_5_28;
wire [31:0] wRegOut_5_28;
wire [31:0] wRegInTop_5_29;
wire [0:0] wRegEnTop_5_29;
wire [31:0] wRegInBot_5_29;
wire [0:0] wRegEnBot_5_29;
wire [31:0] wRegOut_5_29;
wire [31:0] wRegInTop_5_30;
wire [0:0] wRegEnTop_5_30;
wire [31:0] wRegInBot_5_30;
wire [0:0] wRegEnBot_5_30;
wire [31:0] wRegOut_5_30;
wire [31:0] wRegInTop_5_31;
wire [0:0] wRegEnTop_5_31;
wire [31:0] wRegInBot_5_31;
wire [0:0] wRegEnBot_5_31;
wire [31:0] wRegOut_5_31;
wire [0:0] wCtrlOut_6;
wire [0:0] wEnable_6;
wire [31:0] wRegInTop_6_0;
wire [0:0] wRegEnTop_6_0;
wire [31:0] wRegInBot_6_0;
wire [0:0] wRegEnBot_6_0;
wire [31:0] wRegOut_6_0;
wire [31:0] wRegInTop_6_1;
wire [0:0] wRegEnTop_6_1;
wire [31:0] wRegInBot_6_1;
wire [0:0] wRegEnBot_6_1;
wire [31:0] wRegOut_6_1;
wire [31:0] wRegInTop_6_2;
wire [0:0] wRegEnTop_6_2;
wire [31:0] wRegInBot_6_2;
wire [0:0] wRegEnBot_6_2;
wire [31:0] wRegOut_6_2;
wire [31:0] wRegInTop_6_3;
wire [0:0] wRegEnTop_6_3;
wire [31:0] wRegInBot_6_3;
wire [0:0] wRegEnBot_6_3;
wire [31:0] wRegOut_6_3;
wire [31:0] wRegInTop_6_4;
wire [0:0] wRegEnTop_6_4;
wire [31:0] wRegInBot_6_4;
wire [0:0] wRegEnBot_6_4;
wire [31:0] wRegOut_6_4;
wire [31:0] wRegInTop_6_5;
wire [0:0] wRegEnTop_6_5;
wire [31:0] wRegInBot_6_5;
wire [0:0] wRegEnBot_6_5;
wire [31:0] wRegOut_6_5;
wire [31:0] wRegInTop_6_6;
wire [0:0] wRegEnTop_6_6;
wire [31:0] wRegInBot_6_6;
wire [0:0] wRegEnBot_6_6;
wire [31:0] wRegOut_6_6;
wire [31:0] wRegInTop_6_7;
wire [0:0] wRegEnTop_6_7;
wire [31:0] wRegInBot_6_7;
wire [0:0] wRegEnBot_6_7;
wire [31:0] wRegOut_6_7;
wire [31:0] wRegInTop_6_8;
wire [0:0] wRegEnTop_6_8;
wire [31:0] wRegInBot_6_8;
wire [0:0] wRegEnBot_6_8;
wire [31:0] wRegOut_6_8;
wire [31:0] wRegInTop_6_9;
wire [0:0] wRegEnTop_6_9;
wire [31:0] wRegInBot_6_9;
wire [0:0] wRegEnBot_6_9;
wire [31:0] wRegOut_6_9;
wire [31:0] wRegInTop_6_10;
wire [0:0] wRegEnTop_6_10;
wire [31:0] wRegInBot_6_10;
wire [0:0] wRegEnBot_6_10;
wire [31:0] wRegOut_6_10;
wire [31:0] wRegInTop_6_11;
wire [0:0] wRegEnTop_6_11;
wire [31:0] wRegInBot_6_11;
wire [0:0] wRegEnBot_6_11;
wire [31:0] wRegOut_6_11;
wire [31:0] wRegInTop_6_12;
wire [0:0] wRegEnTop_6_12;
wire [31:0] wRegInBot_6_12;
wire [0:0] wRegEnBot_6_12;
wire [31:0] wRegOut_6_12;
wire [31:0] wRegInTop_6_13;
wire [0:0] wRegEnTop_6_13;
wire [31:0] wRegInBot_6_13;
wire [0:0] wRegEnBot_6_13;
wire [31:0] wRegOut_6_13;
wire [31:0] wRegInTop_6_14;
wire [0:0] wRegEnTop_6_14;
wire [31:0] wRegInBot_6_14;
wire [0:0] wRegEnBot_6_14;
wire [31:0] wRegOut_6_14;
wire [31:0] wRegInTop_6_15;
wire [0:0] wRegEnTop_6_15;
wire [31:0] wRegInBot_6_15;
wire [0:0] wRegEnBot_6_15;
wire [31:0] wRegOut_6_15;
wire [31:0] wRegInTop_6_16;
wire [0:0] wRegEnTop_6_16;
wire [31:0] wRegInBot_6_16;
wire [0:0] wRegEnBot_6_16;
wire [31:0] wRegOut_6_16;
wire [31:0] wRegInTop_6_17;
wire [0:0] wRegEnTop_6_17;
wire [31:0] wRegInBot_6_17;
wire [0:0] wRegEnBot_6_17;
wire [31:0] wRegOut_6_17;
wire [31:0] wRegInTop_6_18;
wire [0:0] wRegEnTop_6_18;
wire [31:0] wRegInBot_6_18;
wire [0:0] wRegEnBot_6_18;
wire [31:0] wRegOut_6_18;
wire [31:0] wRegInTop_6_19;
wire [0:0] wRegEnTop_6_19;
wire [31:0] wRegInBot_6_19;
wire [0:0] wRegEnBot_6_19;
wire [31:0] wRegOut_6_19;
wire [31:0] wRegInTop_6_20;
wire [0:0] wRegEnTop_6_20;
wire [31:0] wRegInBot_6_20;
wire [0:0] wRegEnBot_6_20;
wire [31:0] wRegOut_6_20;
wire [31:0] wRegInTop_6_21;
wire [0:0] wRegEnTop_6_21;
wire [31:0] wRegInBot_6_21;
wire [0:0] wRegEnBot_6_21;
wire [31:0] wRegOut_6_21;
wire [31:0] wRegInTop_6_22;
wire [0:0] wRegEnTop_6_22;
wire [31:0] wRegInBot_6_22;
wire [0:0] wRegEnBot_6_22;
wire [31:0] wRegOut_6_22;
wire [31:0] wRegInTop_6_23;
wire [0:0] wRegEnTop_6_23;
wire [31:0] wRegInBot_6_23;
wire [0:0] wRegEnBot_6_23;
wire [31:0] wRegOut_6_23;
wire [31:0] wRegInTop_6_24;
wire [0:0] wRegEnTop_6_24;
wire [31:0] wRegInBot_6_24;
wire [0:0] wRegEnBot_6_24;
wire [31:0] wRegOut_6_24;
wire [31:0] wRegInTop_6_25;
wire [0:0] wRegEnTop_6_25;
wire [31:0] wRegInBot_6_25;
wire [0:0] wRegEnBot_6_25;
wire [31:0] wRegOut_6_25;
wire [31:0] wRegInTop_6_26;
wire [0:0] wRegEnTop_6_26;
wire [31:0] wRegInBot_6_26;
wire [0:0] wRegEnBot_6_26;
wire [31:0] wRegOut_6_26;
wire [31:0] wRegInTop_6_27;
wire [0:0] wRegEnTop_6_27;
wire [31:0] wRegInBot_6_27;
wire [0:0] wRegEnBot_6_27;
wire [31:0] wRegOut_6_27;
wire [31:0] wRegInTop_6_28;
wire [0:0] wRegEnTop_6_28;
wire [31:0] wRegInBot_6_28;
wire [0:0] wRegEnBot_6_28;
wire [31:0] wRegOut_6_28;
wire [31:0] wRegInTop_6_29;
wire [0:0] wRegEnTop_6_29;
wire [31:0] wRegInBot_6_29;
wire [0:0] wRegEnBot_6_29;
wire [31:0] wRegOut_6_29;
wire [31:0] wRegInTop_6_30;
wire [0:0] wRegEnTop_6_30;
wire [31:0] wRegInBot_6_30;
wire [0:0] wRegEnBot_6_30;
wire [31:0] wRegOut_6_30;
wire [31:0] wRegInTop_6_31;
wire [0:0] wRegEnTop_6_31;
wire [31:0] wRegInBot_6_31;
wire [0:0] wRegEnBot_6_31;
wire [31:0] wRegOut_6_31;
wire [31:0] wRegInTop_6_32;
wire [0:0] wRegEnTop_6_32;
wire [31:0] wRegInBot_6_32;
wire [0:0] wRegEnBot_6_32;
wire [31:0] wRegOut_6_32;
wire [31:0] wRegInTop_6_33;
wire [0:0] wRegEnTop_6_33;
wire [31:0] wRegInBot_6_33;
wire [0:0] wRegEnBot_6_33;
wire [31:0] wRegOut_6_33;
wire [31:0] wRegInTop_6_34;
wire [0:0] wRegEnTop_6_34;
wire [31:0] wRegInBot_6_34;
wire [0:0] wRegEnBot_6_34;
wire [31:0] wRegOut_6_34;
wire [31:0] wRegInTop_6_35;
wire [0:0] wRegEnTop_6_35;
wire [31:0] wRegInBot_6_35;
wire [0:0] wRegEnBot_6_35;
wire [31:0] wRegOut_6_35;
wire [31:0] wRegInTop_6_36;
wire [0:0] wRegEnTop_6_36;
wire [31:0] wRegInBot_6_36;
wire [0:0] wRegEnBot_6_36;
wire [31:0] wRegOut_6_36;
wire [31:0] wRegInTop_6_37;
wire [0:0] wRegEnTop_6_37;
wire [31:0] wRegInBot_6_37;
wire [0:0] wRegEnBot_6_37;
wire [31:0] wRegOut_6_37;
wire [31:0] wRegInTop_6_38;
wire [0:0] wRegEnTop_6_38;
wire [31:0] wRegInBot_6_38;
wire [0:0] wRegEnBot_6_38;
wire [31:0] wRegOut_6_38;
wire [31:0] wRegInTop_6_39;
wire [0:0] wRegEnTop_6_39;
wire [31:0] wRegInBot_6_39;
wire [0:0] wRegEnBot_6_39;
wire [31:0] wRegOut_6_39;
wire [31:0] wRegInTop_6_40;
wire [0:0] wRegEnTop_6_40;
wire [31:0] wRegInBot_6_40;
wire [0:0] wRegEnBot_6_40;
wire [31:0] wRegOut_6_40;
wire [31:0] wRegInTop_6_41;
wire [0:0] wRegEnTop_6_41;
wire [31:0] wRegInBot_6_41;
wire [0:0] wRegEnBot_6_41;
wire [31:0] wRegOut_6_41;
wire [31:0] wRegInTop_6_42;
wire [0:0] wRegEnTop_6_42;
wire [31:0] wRegInBot_6_42;
wire [0:0] wRegEnBot_6_42;
wire [31:0] wRegOut_6_42;
wire [31:0] wRegInTop_6_43;
wire [0:0] wRegEnTop_6_43;
wire [31:0] wRegInBot_6_43;
wire [0:0] wRegEnBot_6_43;
wire [31:0] wRegOut_6_43;
wire [31:0] wRegInTop_6_44;
wire [0:0] wRegEnTop_6_44;
wire [31:0] wRegInBot_6_44;
wire [0:0] wRegEnBot_6_44;
wire [31:0] wRegOut_6_44;
wire [31:0] wRegInTop_6_45;
wire [0:0] wRegEnTop_6_45;
wire [31:0] wRegInBot_6_45;
wire [0:0] wRegEnBot_6_45;
wire [31:0] wRegOut_6_45;
wire [31:0] wRegInTop_6_46;
wire [0:0] wRegEnTop_6_46;
wire [31:0] wRegInBot_6_46;
wire [0:0] wRegEnBot_6_46;
wire [31:0] wRegOut_6_46;
wire [31:0] wRegInTop_6_47;
wire [0:0] wRegEnTop_6_47;
wire [31:0] wRegInBot_6_47;
wire [0:0] wRegEnBot_6_47;
wire [31:0] wRegOut_6_47;
wire [31:0] wRegInTop_6_48;
wire [0:0] wRegEnTop_6_48;
wire [31:0] wRegInBot_6_48;
wire [0:0] wRegEnBot_6_48;
wire [31:0] wRegOut_6_48;
wire [31:0] wRegInTop_6_49;
wire [0:0] wRegEnTop_6_49;
wire [31:0] wRegInBot_6_49;
wire [0:0] wRegEnBot_6_49;
wire [31:0] wRegOut_6_49;
wire [31:0] wRegInTop_6_50;
wire [0:0] wRegEnTop_6_50;
wire [31:0] wRegInBot_6_50;
wire [0:0] wRegEnBot_6_50;
wire [31:0] wRegOut_6_50;
wire [31:0] wRegInTop_6_51;
wire [0:0] wRegEnTop_6_51;
wire [31:0] wRegInBot_6_51;
wire [0:0] wRegEnBot_6_51;
wire [31:0] wRegOut_6_51;
wire [31:0] wRegInTop_6_52;
wire [0:0] wRegEnTop_6_52;
wire [31:0] wRegInBot_6_52;
wire [0:0] wRegEnBot_6_52;
wire [31:0] wRegOut_6_52;
wire [31:0] wRegInTop_6_53;
wire [0:0] wRegEnTop_6_53;
wire [31:0] wRegInBot_6_53;
wire [0:0] wRegEnBot_6_53;
wire [31:0] wRegOut_6_53;
wire [31:0] wRegInTop_6_54;
wire [0:0] wRegEnTop_6_54;
wire [31:0] wRegInBot_6_54;
wire [0:0] wRegEnBot_6_54;
wire [31:0] wRegOut_6_54;
wire [31:0] wRegInTop_6_55;
wire [0:0] wRegEnTop_6_55;
wire [31:0] wRegInBot_6_55;
wire [0:0] wRegEnBot_6_55;
wire [31:0] wRegOut_6_55;
wire [31:0] wRegInTop_6_56;
wire [0:0] wRegEnTop_6_56;
wire [31:0] wRegInBot_6_56;
wire [0:0] wRegEnBot_6_56;
wire [31:0] wRegOut_6_56;
wire [31:0] wRegInTop_6_57;
wire [0:0] wRegEnTop_6_57;
wire [31:0] wRegInBot_6_57;
wire [0:0] wRegEnBot_6_57;
wire [31:0] wRegOut_6_57;
wire [31:0] wRegInTop_6_58;
wire [0:0] wRegEnTop_6_58;
wire [31:0] wRegInBot_6_58;
wire [0:0] wRegEnBot_6_58;
wire [31:0] wRegOut_6_58;
wire [31:0] wRegInTop_6_59;
wire [0:0] wRegEnTop_6_59;
wire [31:0] wRegInBot_6_59;
wire [0:0] wRegEnBot_6_59;
wire [31:0] wRegOut_6_59;
wire [31:0] wRegInTop_6_60;
wire [0:0] wRegEnTop_6_60;
wire [31:0] wRegInBot_6_60;
wire [0:0] wRegEnBot_6_60;
wire [31:0] wRegOut_6_60;
wire [31:0] wRegInTop_6_61;
wire [0:0] wRegEnTop_6_61;
wire [31:0] wRegInBot_6_61;
wire [0:0] wRegEnBot_6_61;
wire [31:0] wRegOut_6_61;
wire [31:0] wRegInTop_6_62;
wire [0:0] wRegEnTop_6_62;
wire [31:0] wRegInBot_6_62;
wire [0:0] wRegEnBot_6_62;
wire [31:0] wRegOut_6_62;
wire [31:0] wRegInTop_6_63;
wire [0:0] wRegEnTop_6_63;
wire [31:0] wRegInBot_6_63;
wire [0:0] wRegEnBot_6_63;
wire [31:0] wRegOut_6_63;
wire [0:0] wCtrlOut_7;
wire [0:0] wEnable_7;
wire [31:0] wRegInTop_7_0;
wire [0:0] wRegEnTop_7_0;
wire [31:0] wRegOut_7_0;
wire [31:0] wRegInTop_7_1;
wire [0:0] wRegEnTop_7_1;
wire [31:0] wRegOut_7_1;
wire [31:0] wRegInTop_7_2;
wire [0:0] wRegEnTop_7_2;
wire [31:0] wRegOut_7_2;
wire [31:0] wRegInTop_7_3;
wire [0:0] wRegEnTop_7_3;
wire [31:0] wRegOut_7_3;
wire [31:0] wRegInTop_7_4;
wire [0:0] wRegEnTop_7_4;
wire [31:0] wRegOut_7_4;
wire [31:0] wRegInTop_7_5;
wire [0:0] wRegEnTop_7_5;
wire [31:0] wRegOut_7_5;
wire [31:0] wRegInTop_7_6;
wire [0:0] wRegEnTop_7_6;
wire [31:0] wRegOut_7_6;
wire [31:0] wRegInTop_7_7;
wire [0:0] wRegEnTop_7_7;
wire [31:0] wRegOut_7_7;
wire [31:0] wRegInTop_7_8;
wire [0:0] wRegEnTop_7_8;
wire [31:0] wRegOut_7_8;
wire [31:0] wRegInTop_7_9;
wire [0:0] wRegEnTop_7_9;
wire [31:0] wRegOut_7_9;
wire [31:0] wRegInTop_7_10;
wire [0:0] wRegEnTop_7_10;
wire [31:0] wRegOut_7_10;
wire [31:0] wRegInTop_7_11;
wire [0:0] wRegEnTop_7_11;
wire [31:0] wRegOut_7_11;
wire [31:0] wRegInTop_7_12;
wire [0:0] wRegEnTop_7_12;
wire [31:0] wRegOut_7_12;
wire [31:0] wRegInTop_7_13;
wire [0:0] wRegEnTop_7_13;
wire [31:0] wRegOut_7_13;
wire [31:0] wRegInTop_7_14;
wire [0:0] wRegEnTop_7_14;
wire [31:0] wRegOut_7_14;
wire [31:0] wRegInTop_7_15;
wire [0:0] wRegEnTop_7_15;
wire [31:0] wRegOut_7_15;
wire [31:0] wRegInTop_7_16;
wire [0:0] wRegEnTop_7_16;
wire [31:0] wRegOut_7_16;
wire [31:0] wRegInTop_7_17;
wire [0:0] wRegEnTop_7_17;
wire [31:0] wRegOut_7_17;
wire [31:0] wRegInTop_7_18;
wire [0:0] wRegEnTop_7_18;
wire [31:0] wRegOut_7_18;
wire [31:0] wRegInTop_7_19;
wire [0:0] wRegEnTop_7_19;
wire [31:0] wRegOut_7_19;
wire [31:0] wRegInTop_7_20;
wire [0:0] wRegEnTop_7_20;
wire [31:0] wRegOut_7_20;
wire [31:0] wRegInTop_7_21;
wire [0:0] wRegEnTop_7_21;
wire [31:0] wRegOut_7_21;
wire [31:0] wRegInTop_7_22;
wire [0:0] wRegEnTop_7_22;
wire [31:0] wRegOut_7_22;
wire [31:0] wRegInTop_7_23;
wire [0:0] wRegEnTop_7_23;
wire [31:0] wRegOut_7_23;
wire [31:0] wRegInTop_7_24;
wire [0:0] wRegEnTop_7_24;
wire [31:0] wRegOut_7_24;
wire [31:0] wRegInTop_7_25;
wire [0:0] wRegEnTop_7_25;
wire [31:0] wRegOut_7_25;
wire [31:0] wRegInTop_7_26;
wire [0:0] wRegEnTop_7_26;
wire [31:0] wRegOut_7_26;
wire [31:0] wRegInTop_7_27;
wire [0:0] wRegEnTop_7_27;
wire [31:0] wRegOut_7_27;
wire [31:0] wRegInTop_7_28;
wire [0:0] wRegEnTop_7_28;
wire [31:0] wRegOut_7_28;
wire [31:0] wRegInTop_7_29;
wire [0:0] wRegEnTop_7_29;
wire [31:0] wRegOut_7_29;
wire [31:0] wRegInTop_7_30;
wire [0:0] wRegEnTop_7_30;
wire [31:0] wRegOut_7_30;
wire [31:0] wRegInTop_7_31;
wire [0:0] wRegEnTop_7_31;
wire [31:0] wRegOut_7_31;
wire [31:0] wRegInTop_7_32;
wire [0:0] wRegEnTop_7_32;
wire [31:0] wRegOut_7_32;
wire [31:0] wRegInTop_7_33;
wire [0:0] wRegEnTop_7_33;
wire [31:0] wRegOut_7_33;
wire [31:0] wRegInTop_7_34;
wire [0:0] wRegEnTop_7_34;
wire [31:0] wRegOut_7_34;
wire [31:0] wRegInTop_7_35;
wire [0:0] wRegEnTop_7_35;
wire [31:0] wRegOut_7_35;
wire [31:0] wRegInTop_7_36;
wire [0:0] wRegEnTop_7_36;
wire [31:0] wRegOut_7_36;
wire [31:0] wRegInTop_7_37;
wire [0:0] wRegEnTop_7_37;
wire [31:0] wRegOut_7_37;
wire [31:0] wRegInTop_7_38;
wire [0:0] wRegEnTop_7_38;
wire [31:0] wRegOut_7_38;
wire [31:0] wRegInTop_7_39;
wire [0:0] wRegEnTop_7_39;
wire [31:0] wRegOut_7_39;
wire [31:0] wRegInTop_7_40;
wire [0:0] wRegEnTop_7_40;
wire [31:0] wRegOut_7_40;
wire [31:0] wRegInTop_7_41;
wire [0:0] wRegEnTop_7_41;
wire [31:0] wRegOut_7_41;
wire [31:0] wRegInTop_7_42;
wire [0:0] wRegEnTop_7_42;
wire [31:0] wRegOut_7_42;
wire [31:0] wRegInTop_7_43;
wire [0:0] wRegEnTop_7_43;
wire [31:0] wRegOut_7_43;
wire [31:0] wRegInTop_7_44;
wire [0:0] wRegEnTop_7_44;
wire [31:0] wRegOut_7_44;
wire [31:0] wRegInTop_7_45;
wire [0:0] wRegEnTop_7_45;
wire [31:0] wRegOut_7_45;
wire [31:0] wRegInTop_7_46;
wire [0:0] wRegEnTop_7_46;
wire [31:0] wRegOut_7_46;
wire [31:0] wRegInTop_7_47;
wire [0:0] wRegEnTop_7_47;
wire [31:0] wRegOut_7_47;
wire [31:0] wRegInTop_7_48;
wire [0:0] wRegEnTop_7_48;
wire [31:0] wRegOut_7_48;
wire [31:0] wRegInTop_7_49;
wire [0:0] wRegEnTop_7_49;
wire [31:0] wRegOut_7_49;
wire [31:0] wRegInTop_7_50;
wire [0:0] wRegEnTop_7_50;
wire [31:0] wRegOut_7_50;
wire [31:0] wRegInTop_7_51;
wire [0:0] wRegEnTop_7_51;
wire [31:0] wRegOut_7_51;
wire [31:0] wRegInTop_7_52;
wire [0:0] wRegEnTop_7_52;
wire [31:0] wRegOut_7_52;
wire [31:0] wRegInTop_7_53;
wire [0:0] wRegEnTop_7_53;
wire [31:0] wRegOut_7_53;
wire [31:0] wRegInTop_7_54;
wire [0:0] wRegEnTop_7_54;
wire [31:0] wRegOut_7_54;
wire [31:0] wRegInTop_7_55;
wire [0:0] wRegEnTop_7_55;
wire [31:0] wRegOut_7_55;
wire [31:0] wRegInTop_7_56;
wire [0:0] wRegEnTop_7_56;
wire [31:0] wRegOut_7_56;
wire [31:0] wRegInTop_7_57;
wire [0:0] wRegEnTop_7_57;
wire [31:0] wRegOut_7_57;
wire [31:0] wRegInTop_7_58;
wire [0:0] wRegEnTop_7_58;
wire [31:0] wRegOut_7_58;
wire [31:0] wRegInTop_7_59;
wire [0:0] wRegEnTop_7_59;
wire [31:0] wRegOut_7_59;
wire [31:0] wRegInTop_7_60;
wire [0:0] wRegEnTop_7_60;
wire [31:0] wRegOut_7_60;
wire [31:0] wRegInTop_7_61;
wire [0:0] wRegEnTop_7_61;
wire [31:0] wRegOut_7_61;
wire [31:0] wRegInTop_7_62;
wire [0:0] wRegEnTop_7_62;
wire [31:0] wRegOut_7_62;
wire [31:0] wRegInTop_7_63;
wire [0:0] wRegEnTop_7_63;
wire [31:0] wRegOut_7_63;
wire [31:0] wRegInTop_7_64;
wire [0:0] wRegEnTop_7_64;
wire [31:0] wRegOut_7_64;
wire [31:0] wRegInTop_7_65;
wire [0:0] wRegEnTop_7_65;
wire [31:0] wRegOut_7_65;
wire [31:0] wRegInTop_7_66;
wire [0:0] wRegEnTop_7_66;
wire [31:0] wRegOut_7_66;
wire [31:0] wRegInTop_7_67;
wire [0:0] wRegEnTop_7_67;
wire [31:0] wRegOut_7_67;
wire [31:0] wRegInTop_7_68;
wire [0:0] wRegEnTop_7_68;
wire [31:0] wRegOut_7_68;
wire [31:0] wRegInTop_7_69;
wire [0:0] wRegEnTop_7_69;
wire [31:0] wRegOut_7_69;
wire [31:0] wRegInTop_7_70;
wire [0:0] wRegEnTop_7_70;
wire [31:0] wRegOut_7_70;
wire [31:0] wRegInTop_7_71;
wire [0:0] wRegEnTop_7_71;
wire [31:0] wRegOut_7_71;
wire [31:0] wRegInTop_7_72;
wire [0:0] wRegEnTop_7_72;
wire [31:0] wRegOut_7_72;
wire [31:0] wRegInTop_7_73;
wire [0:0] wRegEnTop_7_73;
wire [31:0] wRegOut_7_73;
wire [31:0] wRegInTop_7_74;
wire [0:0] wRegEnTop_7_74;
wire [31:0] wRegOut_7_74;
wire [31:0] wRegInTop_7_75;
wire [0:0] wRegEnTop_7_75;
wire [31:0] wRegOut_7_75;
wire [31:0] wRegInTop_7_76;
wire [0:0] wRegEnTop_7_76;
wire [31:0] wRegOut_7_76;
wire [31:0] wRegInTop_7_77;
wire [0:0] wRegEnTop_7_77;
wire [31:0] wRegOut_7_77;
wire [31:0] wRegInTop_7_78;
wire [0:0] wRegEnTop_7_78;
wire [31:0] wRegOut_7_78;
wire [31:0] wRegInTop_7_79;
wire [0:0] wRegEnTop_7_79;
wire [31:0] wRegOut_7_79;
wire [31:0] wRegInTop_7_80;
wire [0:0] wRegEnTop_7_80;
wire [31:0] wRegOut_7_80;
wire [31:0] wRegInTop_7_81;
wire [0:0] wRegEnTop_7_81;
wire [31:0] wRegOut_7_81;
wire [31:0] wRegInTop_7_82;
wire [0:0] wRegEnTop_7_82;
wire [31:0] wRegOut_7_82;
wire [31:0] wRegInTop_7_83;
wire [0:0] wRegEnTop_7_83;
wire [31:0] wRegOut_7_83;
wire [31:0] wRegInTop_7_84;
wire [0:0] wRegEnTop_7_84;
wire [31:0] wRegOut_7_84;
wire [31:0] wRegInTop_7_85;
wire [0:0] wRegEnTop_7_85;
wire [31:0] wRegOut_7_85;
wire [31:0] wRegInTop_7_86;
wire [0:0] wRegEnTop_7_86;
wire [31:0] wRegOut_7_86;
wire [31:0] wRegInTop_7_87;
wire [0:0] wRegEnTop_7_87;
wire [31:0] wRegOut_7_87;
wire [31:0] wRegInTop_7_88;
wire [0:0] wRegEnTop_7_88;
wire [31:0] wRegOut_7_88;
wire [31:0] wRegInTop_7_89;
wire [0:0] wRegEnTop_7_89;
wire [31:0] wRegOut_7_89;
wire [31:0] wRegInTop_7_90;
wire [0:0] wRegEnTop_7_90;
wire [31:0] wRegOut_7_90;
wire [31:0] wRegInTop_7_91;
wire [0:0] wRegEnTop_7_91;
wire [31:0] wRegOut_7_91;
wire [31:0] wRegInTop_7_92;
wire [0:0] wRegEnTop_7_92;
wire [31:0] wRegOut_7_92;
wire [31:0] wRegInTop_7_93;
wire [0:0] wRegEnTop_7_93;
wire [31:0] wRegOut_7_93;
wire [31:0] wRegInTop_7_94;
wire [0:0] wRegEnTop_7_94;
wire [31:0] wRegOut_7_94;
wire [31:0] wRegInTop_7_95;
wire [0:0] wRegEnTop_7_95;
wire [31:0] wRegOut_7_95;
wire [31:0] wRegInTop_7_96;
wire [0:0] wRegEnTop_7_96;
wire [31:0] wRegOut_7_96;
wire [31:0] wRegInTop_7_97;
wire [0:0] wRegEnTop_7_97;
wire [31:0] wRegOut_7_97;
wire [31:0] wRegInTop_7_98;
wire [0:0] wRegEnTop_7_98;
wire [31:0] wRegOut_7_98;
wire [31:0] wRegInTop_7_99;
wire [0:0] wRegEnTop_7_99;
wire [31:0] wRegOut_7_99;
wire [31:0] wRegInTop_7_100;
wire [0:0] wRegEnTop_7_100;
wire [31:0] wRegOut_7_100;
wire [31:0] wRegInTop_7_101;
wire [0:0] wRegEnTop_7_101;
wire [31:0] wRegOut_7_101;
wire [31:0] wRegInTop_7_102;
wire [0:0] wRegEnTop_7_102;
wire [31:0] wRegOut_7_102;
wire [31:0] wRegInTop_7_103;
wire [0:0] wRegEnTop_7_103;
wire [31:0] wRegOut_7_103;
wire [31:0] wRegInTop_7_104;
wire [0:0] wRegEnTop_7_104;
wire [31:0] wRegOut_7_104;
wire [31:0] wRegInTop_7_105;
wire [0:0] wRegEnTop_7_105;
wire [31:0] wRegOut_7_105;
wire [31:0] wRegInTop_7_106;
wire [0:0] wRegEnTop_7_106;
wire [31:0] wRegOut_7_106;
wire [31:0] wRegInTop_7_107;
wire [0:0] wRegEnTop_7_107;
wire [31:0] wRegOut_7_107;
wire [31:0] wRegInTop_7_108;
wire [0:0] wRegEnTop_7_108;
wire [31:0] wRegOut_7_108;
wire [31:0] wRegInTop_7_109;
wire [0:0] wRegEnTop_7_109;
wire [31:0] wRegOut_7_109;
wire [31:0] wRegInTop_7_110;
wire [0:0] wRegEnTop_7_110;
wire [31:0] wRegOut_7_110;
wire [31:0] wRegInTop_7_111;
wire [0:0] wRegEnTop_7_111;
wire [31:0] wRegOut_7_111;
wire [31:0] wRegInTop_7_112;
wire [0:0] wRegEnTop_7_112;
wire [31:0] wRegOut_7_112;
wire [31:0] wRegInTop_7_113;
wire [0:0] wRegEnTop_7_113;
wire [31:0] wRegOut_7_113;
wire [31:0] wRegInTop_7_114;
wire [0:0] wRegEnTop_7_114;
wire [31:0] wRegOut_7_114;
wire [31:0] wRegInTop_7_115;
wire [0:0] wRegEnTop_7_115;
wire [31:0] wRegOut_7_115;
wire [31:0] wRegInTop_7_116;
wire [0:0] wRegEnTop_7_116;
wire [31:0] wRegOut_7_116;
wire [31:0] wRegInTop_7_117;
wire [0:0] wRegEnTop_7_117;
wire [31:0] wRegOut_7_117;
wire [31:0] wRegInTop_7_118;
wire [0:0] wRegEnTop_7_118;
wire [31:0] wRegOut_7_118;
wire [31:0] wRegInTop_7_119;
wire [0:0] wRegEnTop_7_119;
wire [31:0] wRegOut_7_119;
wire [31:0] wRegInTop_7_120;
wire [0:0] wRegEnTop_7_120;
wire [31:0] wRegOut_7_120;
wire [31:0] wRegInTop_7_121;
wire [0:0] wRegEnTop_7_121;
wire [31:0] wRegOut_7_121;
wire [31:0] wRegInTop_7_122;
wire [0:0] wRegEnTop_7_122;
wire [31:0] wRegOut_7_122;
wire [31:0] wRegInTop_7_123;
wire [0:0] wRegEnTop_7_123;
wire [31:0] wRegOut_7_123;
wire [31:0] wRegInTop_7_124;
wire [0:0] wRegEnTop_7_124;
wire [31:0] wRegOut_7_124;
wire [31:0] wRegInTop_7_125;
wire [0:0] wRegEnTop_7_125;
wire [31:0] wRegOut_7_125;
wire [31:0] wRegInTop_7_126;
wire [0:0] wRegEnTop_7_126;
wire [31:0] wRegOut_7_126;
wire [31:0] wRegInTop_7_127;
wire [0:0] wRegEnTop_7_127;
wire [31:0] wRegOut_7_127;
wire [0:0] ScanEnable;
wire [31:0] ScanLink0;
wire [31:0] ScanLink1;
wire [31:0] ScanLink2;
wire [31:0] ScanLink3;
wire [31:0] ScanLink4;
wire [31:0] ScanLink5;
wire [31:0] ScanLink6;
wire [31:0] ScanLink7;
wire [31:0] ScanLink8;
wire [31:0] ScanLink9;
wire [31:0] ScanLink10;
wire [31:0] ScanLink11;
wire [31:0] ScanLink12;
wire [31:0] ScanLink13;
wire [31:0] ScanLink14;
wire [31:0] ScanLink15;
wire [31:0] ScanLink16;
wire [31:0] ScanLink17;
wire [31:0] ScanLink18;
wire [31:0] ScanLink19;
wire [31:0] ScanLink20;
wire [31:0] ScanLink21;
wire [31:0] ScanLink22;
wire [31:0] ScanLink23;
wire [31:0] ScanLink24;
wire [31:0] ScanLink25;
wire [31:0] ScanLink26;
wire [31:0] ScanLink27;
wire [31:0] ScanLink28;
wire [31:0] ScanLink29;
wire [31:0] ScanLink30;
wire [31:0] ScanLink31;
wire [31:0] ScanLink32;
wire [31:0] ScanLink33;
wire [31:0] ScanLink34;
wire [31:0] ScanLink35;
wire [31:0] ScanLink36;
wire [31:0] ScanLink37;
wire [31:0] ScanLink38;
wire [31:0] ScanLink39;
wire [31:0] ScanLink40;
wire [31:0] ScanLink41;
wire [31:0] ScanLink42;
wire [31:0] ScanLink43;
wire [31:0] ScanLink44;
wire [31:0] ScanLink45;
wire [31:0] ScanLink46;
wire [31:0] ScanLink47;
wire [31:0] ScanLink48;
wire [31:0] ScanLink49;
wire [31:0] ScanLink50;
wire [31:0] ScanLink51;
wire [31:0] ScanLink52;
wire [31:0] ScanLink53;
wire [31:0] ScanLink54;
wire [31:0] ScanLink55;
wire [31:0] ScanLink56;
wire [31:0] ScanLink57;
wire [31:0] ScanLink58;
wire [31:0] ScanLink59;
wire [31:0] ScanLink60;
wire [31:0] ScanLink61;
wire [31:0] ScanLink62;
wire [31:0] ScanLink63;
wire [31:0] ScanLink64;
wire [31:0] ScanLink65;
wire [31:0] ScanLink66;
wire [31:0] ScanLink67;
wire [31:0] ScanLink68;
wire [31:0] ScanLink69;
wire [31:0] ScanLink70;
wire [31:0] ScanLink71;
wire [31:0] ScanLink72;
wire [31:0] ScanLink73;
wire [31:0] ScanLink74;
wire [31:0] ScanLink75;
wire [31:0] ScanLink76;
wire [31:0] ScanLink77;
wire [31:0] ScanLink78;
wire [31:0] ScanLink79;
wire [31:0] ScanLink80;
wire [31:0] ScanLink81;
wire [31:0] ScanLink82;
wire [31:0] ScanLink83;
wire [31:0] ScanLink84;
wire [31:0] ScanLink85;
wire [31:0] ScanLink86;
wire [31:0] ScanLink87;
wire [31:0] ScanLink88;
wire [31:0] ScanLink89;
wire [31:0] ScanLink90;
wire [31:0] ScanLink91;
wire [31:0] ScanLink92;
wire [31:0] ScanLink93;
wire [31:0] ScanLink94;
wire [31:0] ScanLink95;
wire [31:0] ScanLink96;
wire [31:0] ScanLink97;
wire [31:0] ScanLink98;
wire [31:0] ScanLink99;
wire [31:0] ScanLink100;
wire [31:0] ScanLink101;
wire [31:0] ScanLink102;
wire [31:0] ScanLink103;
wire [31:0] ScanLink104;
wire [31:0] ScanLink105;
wire [31:0] ScanLink106;
wire [31:0] ScanLink107;
wire [31:0] ScanLink108;
wire [31:0] ScanLink109;
wire [31:0] ScanLink110;
wire [31:0] ScanLink111;
wire [31:0] ScanLink112;
wire [31:0] ScanLink113;
wire [31:0] ScanLink114;
wire [31:0] ScanLink115;
wire [31:0] ScanLink116;
wire [31:0] ScanLink117;
wire [31:0] ScanLink118;
wire [31:0] ScanLink119;
wire [31:0] ScanLink120;
wire [31:0] ScanLink121;
wire [31:0] ScanLink122;
wire [31:0] ScanLink123;
wire [31:0] ScanLink124;
wire [31:0] ScanLink125;
wire [31:0] ScanLink126;
wire [31:0] ScanLink127;
wire [31:0] ScanLink128;
wire [31:0] ScanLink129;
wire [31:0] ScanLink130;
wire [31:0] ScanLink131;
wire [31:0] ScanLink132;
wire [31:0] ScanLink133;
wire [31:0] ScanLink134;
wire [31:0] ScanLink135;
wire [31:0] ScanLink136;
wire [31:0] ScanLink137;
wire [31:0] ScanLink138;
wire [31:0] ScanLink139;
wire [31:0] ScanLink140;
wire [31:0] ScanLink141;
wire [31:0] ScanLink142;
wire [31:0] ScanLink143;
wire [31:0] ScanLink144;
wire [31:0] ScanLink145;
wire [31:0] ScanLink146;
wire [31:0] ScanLink147;
wire [31:0] ScanLink148;
wire [31:0] ScanLink149;
wire [31:0] ScanLink150;
wire [31:0] ScanLink151;
wire [31:0] ScanLink152;
wire [31:0] ScanLink153;
wire [31:0] ScanLink154;
wire [31:0] ScanLink155;
wire [31:0] ScanLink156;
wire [31:0] ScanLink157;
wire [31:0] ScanLink158;
wire [31:0] ScanLink159;
wire [31:0] ScanLink160;
wire [31:0] ScanLink161;
wire [31:0] ScanLink162;
wire [31:0] ScanLink163;
wire [31:0] ScanLink164;
wire [31:0] ScanLink165;
wire [31:0] ScanLink166;
wire [31:0] ScanLink167;
wire [31:0] ScanLink168;
wire [31:0] ScanLink169;
wire [31:0] ScanLink170;
wire [31:0] ScanLink171;
wire [31:0] ScanLink172;
wire [31:0] ScanLink173;
wire [31:0] ScanLink174;
wire [31:0] ScanLink175;
wire [31:0] ScanLink176;
wire [31:0] ScanLink177;
wire [31:0] ScanLink178;
wire [31:0] ScanLink179;
wire [31:0] ScanLink180;
wire [31:0] ScanLink181;
wire [31:0] ScanLink182;
wire [31:0] ScanLink183;
wire [31:0] ScanLink184;
wire [31:0] ScanLink185;
wire [31:0] ScanLink186;
wire [31:0] ScanLink187;
wire [31:0] ScanLink188;
wire [31:0] ScanLink189;
wire [31:0] ScanLink190;
wire [31:0] ScanLink191;
wire [31:0] ScanLink192;
wire [31:0] ScanLink193;
wire [31:0] ScanLink194;
wire [31:0] ScanLink195;
wire [31:0] ScanLink196;
wire [31:0] ScanLink197;
wire [31:0] ScanLink198;
wire [31:0] ScanLink199;
wire [31:0] ScanLink200;
wire [31:0] ScanLink201;
wire [31:0] ScanLink202;
wire [31:0] ScanLink203;
wire [31:0] ScanLink204;
wire [31:0] ScanLink205;
wire [31:0] ScanLink206;
wire [31:0] ScanLink207;
wire [31:0] ScanLink208;
wire [31:0] ScanLink209;
wire [31:0] ScanLink210;
wire [31:0] ScanLink211;
wire [31:0] ScanLink212;
wire [31:0] ScanLink213;
wire [31:0] ScanLink214;
wire [31:0] ScanLink215;
wire [31:0] ScanLink216;
wire [31:0] ScanLink217;
wire [31:0] ScanLink218;
wire [31:0] ScanLink219;
wire [31:0] ScanLink220;
wire [31:0] ScanLink221;
wire [31:0] ScanLink222;
wire [31:0] ScanLink223;
wire [31:0] ScanLink224;
wire [31:0] ScanLink225;
wire [31:0] ScanLink226;
wire [31:0] ScanLink227;
wire [31:0] ScanLink228;
wire [31:0] ScanLink229;
wire [31:0] ScanLink230;
wire [31:0] ScanLink231;
wire [31:0] ScanLink232;
wire [31:0] ScanLink233;
wire [31:0] ScanLink234;
wire [31:0] ScanLink235;
wire [31:0] ScanLink236;
wire [31:0] ScanLink237;
wire [31:0] ScanLink238;
wire [31:0] ScanLink239;
wire [31:0] ScanLink240;
wire [31:0] ScanLink241;
wire [31:0] ScanLink242;
wire [31:0] ScanLink243;
wire [31:0] ScanLink244;
wire [31:0] ScanLink245;
wire [31:0] ScanLink246;
wire [31:0] ScanLink247;
wire [31:0] ScanLink248;
wire [31:0] ScanLink249;
wire [31:0] ScanLink250;
wire [31:0] ScanLink251;
wire [31:0] ScanLink252;
wire [31:0] ScanLink253;
wire [31:0] ScanLink254;
wire [31:0] ScanLink255;
BHeap_Reg #( 32, 1, 1 ) BHR_0_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_0_0), .Enable1(1'b0), .In1(32'b0), .Enable2(wRegEnBot_0_0), .In2(wRegInBot_0_0), .ScanIn(ScanLink1), .ScanOut(ScanLink0), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_1_0), .Enable1(wRegEnTop_1_0), .In1(wRegInTop_1_0), .Enable2(wRegEnBot_1_0), .In2(wRegInBot_1_0), .ScanIn(ScanLink2), .ScanOut(ScanLink1), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_1_1), .Enable1(wRegEnTop_1_1), .In1(wRegInTop_1_1), .Enable2(wRegEnBot_1_1), .In2(wRegInBot_1_1), .ScanIn(ScanLink3), .ScanOut(ScanLink2), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_2_0), .Enable1(wRegEnTop_2_0), .In1(wRegInTop_2_0), .Enable2(wRegEnBot_2_0), .In2(wRegInBot_2_0), .ScanIn(ScanLink4), .ScanOut(ScanLink3), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_2_1), .Enable1(wRegEnTop_2_1), .In1(wRegInTop_2_1), .Enable2(wRegEnBot_2_1), .In2(wRegInBot_2_1), .ScanIn(ScanLink5), .ScanOut(ScanLink4), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_2_2), .Enable1(wRegEnTop_2_2), .In1(wRegInTop_2_2), .Enable2(wRegEnBot_2_2), .In2(wRegInBot_2_2), .ScanIn(ScanLink6), .ScanOut(ScanLink5), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_2_3), .Enable1(wRegEnTop_2_3), .In1(wRegInTop_2_3), .Enable2(wRegEnBot_2_3), .In2(wRegInBot_2_3), .ScanIn(ScanLink7), .ScanOut(ScanLink6), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_0), .Enable1(wRegEnTop_3_0), .In1(wRegInTop_3_0), .Enable2(wRegEnBot_3_0), .In2(wRegInBot_3_0), .ScanIn(ScanLink8), .ScanOut(ScanLink7), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_1), .Enable1(wRegEnTop_3_1), .In1(wRegInTop_3_1), .Enable2(wRegEnBot_3_1), .In2(wRegInBot_3_1), .ScanIn(ScanLink9), .ScanOut(ScanLink8), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_2), .Enable1(wRegEnTop_3_2), .In1(wRegInTop_3_2), .Enable2(wRegEnBot_3_2), .In2(wRegInBot_3_2), .ScanIn(ScanLink10), .ScanOut(ScanLink9), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_3), .Enable1(wRegEnTop_3_3), .In1(wRegInTop_3_3), .Enable2(wRegEnBot_3_3), .In2(wRegInBot_3_3), .ScanIn(ScanLink11), .ScanOut(ScanLink10), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_4), .Enable1(wRegEnTop_3_4), .In1(wRegInTop_3_4), .Enable2(wRegEnBot_3_4), .In2(wRegInBot_3_4), .ScanIn(ScanLink12), .ScanOut(ScanLink11), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_5), .Enable1(wRegEnTop_3_5), .In1(wRegInTop_3_5), .Enable2(wRegEnBot_3_5), .In2(wRegInBot_3_5), .ScanIn(ScanLink13), .ScanOut(ScanLink12), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_6), .Enable1(wRegEnTop_3_6), .In1(wRegInTop_3_6), .Enable2(wRegEnBot_3_6), .In2(wRegInBot_3_6), .ScanIn(ScanLink14), .ScanOut(ScanLink13), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_3_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_3_7), .Enable1(wRegEnTop_3_7), .In1(wRegInTop_3_7), .Enable2(wRegEnBot_3_7), .In2(wRegInBot_3_7), .ScanIn(ScanLink15), .ScanOut(ScanLink14), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_0), .Enable1(wRegEnTop_4_0), .In1(wRegInTop_4_0), .Enable2(wRegEnBot_4_0), .In2(wRegInBot_4_0), .ScanIn(ScanLink16), .ScanOut(ScanLink15), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_1), .Enable1(wRegEnTop_4_1), .In1(wRegInTop_4_1), .Enable2(wRegEnBot_4_1), .In2(wRegInBot_4_1), .ScanIn(ScanLink17), .ScanOut(ScanLink16), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_2), .Enable1(wRegEnTop_4_2), .In1(wRegInTop_4_2), .Enable2(wRegEnBot_4_2), .In2(wRegInBot_4_2), .ScanIn(ScanLink18), .ScanOut(ScanLink17), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_3), .Enable1(wRegEnTop_4_3), .In1(wRegInTop_4_3), .Enable2(wRegEnBot_4_3), .In2(wRegInBot_4_3), .ScanIn(ScanLink19), .ScanOut(ScanLink18), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_4), .Enable1(wRegEnTop_4_4), .In1(wRegInTop_4_4), .Enable2(wRegEnBot_4_4), .In2(wRegInBot_4_4), .ScanIn(ScanLink20), .ScanOut(ScanLink19), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_5), .Enable1(wRegEnTop_4_5), .In1(wRegInTop_4_5), .Enable2(wRegEnBot_4_5), .In2(wRegInBot_4_5), .ScanIn(ScanLink21), .ScanOut(ScanLink20), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_6), .Enable1(wRegEnTop_4_6), .In1(wRegInTop_4_6), .Enable2(wRegEnBot_4_6), .In2(wRegInBot_4_6), .ScanIn(ScanLink22), .ScanOut(ScanLink21), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_7), .Enable1(wRegEnTop_4_7), .In1(wRegInTop_4_7), .Enable2(wRegEnBot_4_7), .In2(wRegInBot_4_7), .ScanIn(ScanLink23), .ScanOut(ScanLink22), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_8), .Enable1(wRegEnTop_4_8), .In1(wRegInTop_4_8), .Enable2(wRegEnBot_4_8), .In2(wRegInBot_4_8), .ScanIn(ScanLink24), .ScanOut(ScanLink23), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_9), .Enable1(wRegEnTop_4_9), .In1(wRegInTop_4_9), .Enable2(wRegEnBot_4_9), .In2(wRegInBot_4_9), .ScanIn(ScanLink25), .ScanOut(ScanLink24), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_10), .Enable1(wRegEnTop_4_10), .In1(wRegInTop_4_10), .Enable2(wRegEnBot_4_10), .In2(wRegInBot_4_10), .ScanIn(ScanLink26), .ScanOut(ScanLink25), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_11), .Enable1(wRegEnTop_4_11), .In1(wRegInTop_4_11), .Enable2(wRegEnBot_4_11), .In2(wRegInBot_4_11), .ScanIn(ScanLink27), .ScanOut(ScanLink26), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_12), .Enable1(wRegEnTop_4_12), .In1(wRegInTop_4_12), .Enable2(wRegEnBot_4_12), .In2(wRegInBot_4_12), .ScanIn(ScanLink28), .ScanOut(ScanLink27), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_13), .Enable1(wRegEnTop_4_13), .In1(wRegInTop_4_13), .Enable2(wRegEnBot_4_13), .In2(wRegInBot_4_13), .ScanIn(ScanLink29), .ScanOut(ScanLink28), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_14), .Enable1(wRegEnTop_4_14), .In1(wRegInTop_4_14), .Enable2(wRegEnBot_4_14), .In2(wRegInBot_4_14), .ScanIn(ScanLink30), .ScanOut(ScanLink29), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_4_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_4_15), .Enable1(wRegEnTop_4_15), .In1(wRegInTop_4_15), .Enable2(wRegEnBot_4_15), .In2(wRegInBot_4_15), .ScanIn(ScanLink31), .ScanOut(ScanLink30), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_0), .Enable1(wRegEnTop_5_0), .In1(wRegInTop_5_0), .Enable2(wRegEnBot_5_0), .In2(wRegInBot_5_0), .ScanIn(ScanLink32), .ScanOut(ScanLink31), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_1), .Enable1(wRegEnTop_5_1), .In1(wRegInTop_5_1), .Enable2(wRegEnBot_5_1), .In2(wRegInBot_5_1), .ScanIn(ScanLink33), .ScanOut(ScanLink32), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_2), .Enable1(wRegEnTop_5_2), .In1(wRegInTop_5_2), .Enable2(wRegEnBot_5_2), .In2(wRegInBot_5_2), .ScanIn(ScanLink34), .ScanOut(ScanLink33), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_3), .Enable1(wRegEnTop_5_3), .In1(wRegInTop_5_3), .Enable2(wRegEnBot_5_3), .In2(wRegInBot_5_3), .ScanIn(ScanLink35), .ScanOut(ScanLink34), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_4), .Enable1(wRegEnTop_5_4), .In1(wRegInTop_5_4), .Enable2(wRegEnBot_5_4), .In2(wRegInBot_5_4), .ScanIn(ScanLink36), .ScanOut(ScanLink35), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_5), .Enable1(wRegEnTop_5_5), .In1(wRegInTop_5_5), .Enable2(wRegEnBot_5_5), .In2(wRegInBot_5_5), .ScanIn(ScanLink37), .ScanOut(ScanLink36), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_6), .Enable1(wRegEnTop_5_6), .In1(wRegInTop_5_6), .Enable2(wRegEnBot_5_6), .In2(wRegInBot_5_6), .ScanIn(ScanLink38), .ScanOut(ScanLink37), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_7), .Enable1(wRegEnTop_5_7), .In1(wRegInTop_5_7), .Enable2(wRegEnBot_5_7), .In2(wRegInBot_5_7), .ScanIn(ScanLink39), .ScanOut(ScanLink38), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_8), .Enable1(wRegEnTop_5_8), .In1(wRegInTop_5_8), .Enable2(wRegEnBot_5_8), .In2(wRegInBot_5_8), .ScanIn(ScanLink40), .ScanOut(ScanLink39), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_9), .Enable1(wRegEnTop_5_9), .In1(wRegInTop_5_9), .Enable2(wRegEnBot_5_9), .In2(wRegInBot_5_9), .ScanIn(ScanLink41), .ScanOut(ScanLink40), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_10), .Enable1(wRegEnTop_5_10), .In1(wRegInTop_5_10), .Enable2(wRegEnBot_5_10), .In2(wRegInBot_5_10), .ScanIn(ScanLink42), .ScanOut(ScanLink41), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_11), .Enable1(wRegEnTop_5_11), .In1(wRegInTop_5_11), .Enable2(wRegEnBot_5_11), .In2(wRegInBot_5_11), .ScanIn(ScanLink43), .ScanOut(ScanLink42), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_12), .Enable1(wRegEnTop_5_12), .In1(wRegInTop_5_12), .Enable2(wRegEnBot_5_12), .In2(wRegInBot_5_12), .ScanIn(ScanLink44), .ScanOut(ScanLink43), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_13), .Enable1(wRegEnTop_5_13), .In1(wRegInTop_5_13), .Enable2(wRegEnBot_5_13), .In2(wRegInBot_5_13), .ScanIn(ScanLink45), .ScanOut(ScanLink44), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_14), .Enable1(wRegEnTop_5_14), .In1(wRegInTop_5_14), .Enable2(wRegEnBot_5_14), .In2(wRegInBot_5_14), .ScanIn(ScanLink46), .ScanOut(ScanLink45), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_15), .Enable1(wRegEnTop_5_15), .In1(wRegInTop_5_15), .Enable2(wRegEnBot_5_15), .In2(wRegInBot_5_15), .ScanIn(ScanLink47), .ScanOut(ScanLink46), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_16), .Enable1(wRegEnTop_5_16), .In1(wRegInTop_5_16), .Enable2(wRegEnBot_5_16), .In2(wRegInBot_5_16), .ScanIn(ScanLink48), .ScanOut(ScanLink47), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_17), .Enable1(wRegEnTop_5_17), .In1(wRegInTop_5_17), .Enable2(wRegEnBot_5_17), .In2(wRegInBot_5_17), .ScanIn(ScanLink49), .ScanOut(ScanLink48), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_18), .Enable1(wRegEnTop_5_18), .In1(wRegInTop_5_18), .Enable2(wRegEnBot_5_18), .In2(wRegInBot_5_18), .ScanIn(ScanLink50), .ScanOut(ScanLink49), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_19), .Enable1(wRegEnTop_5_19), .In1(wRegInTop_5_19), .Enable2(wRegEnBot_5_19), .In2(wRegInBot_5_19), .ScanIn(ScanLink51), .ScanOut(ScanLink50), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_20), .Enable1(wRegEnTop_5_20), .In1(wRegInTop_5_20), .Enable2(wRegEnBot_5_20), .In2(wRegInBot_5_20), .ScanIn(ScanLink52), .ScanOut(ScanLink51), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_21), .Enable1(wRegEnTop_5_21), .In1(wRegInTop_5_21), .Enable2(wRegEnBot_5_21), .In2(wRegInBot_5_21), .ScanIn(ScanLink53), .ScanOut(ScanLink52), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_22), .Enable1(wRegEnTop_5_22), .In1(wRegInTop_5_22), .Enable2(wRegEnBot_5_22), .In2(wRegInBot_5_22), .ScanIn(ScanLink54), .ScanOut(ScanLink53), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_23), .Enable1(wRegEnTop_5_23), .In1(wRegInTop_5_23), .Enable2(wRegEnBot_5_23), .In2(wRegInBot_5_23), .ScanIn(ScanLink55), .ScanOut(ScanLink54), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_24), .Enable1(wRegEnTop_5_24), .In1(wRegInTop_5_24), .Enable2(wRegEnBot_5_24), .In2(wRegInBot_5_24), .ScanIn(ScanLink56), .ScanOut(ScanLink55), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_25), .Enable1(wRegEnTop_5_25), .In1(wRegInTop_5_25), .Enable2(wRegEnBot_5_25), .In2(wRegInBot_5_25), .ScanIn(ScanLink57), .ScanOut(ScanLink56), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_26), .Enable1(wRegEnTop_5_26), .In1(wRegInTop_5_26), .Enable2(wRegEnBot_5_26), .In2(wRegInBot_5_26), .ScanIn(ScanLink58), .ScanOut(ScanLink57), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_27), .Enable1(wRegEnTop_5_27), .In1(wRegInTop_5_27), .Enable2(wRegEnBot_5_27), .In2(wRegInBot_5_27), .ScanIn(ScanLink59), .ScanOut(ScanLink58), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_28), .Enable1(wRegEnTop_5_28), .In1(wRegInTop_5_28), .Enable2(wRegEnBot_5_28), .In2(wRegInBot_5_28), .ScanIn(ScanLink60), .ScanOut(ScanLink59), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_29), .Enable1(wRegEnTop_5_29), .In1(wRegInTop_5_29), .Enable2(wRegEnBot_5_29), .In2(wRegInBot_5_29), .ScanIn(ScanLink61), .ScanOut(ScanLink60), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_30), .Enable1(wRegEnTop_5_30), .In1(wRegInTop_5_30), .Enable2(wRegEnBot_5_30), .In2(wRegInBot_5_30), .ScanIn(ScanLink62), .ScanOut(ScanLink61), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_5_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_5_31), .Enable1(wRegEnTop_5_31), .In1(wRegInTop_5_31), .Enable2(wRegEnBot_5_31), .In2(wRegInBot_5_31), .ScanIn(ScanLink63), .ScanOut(ScanLink62), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_0), .Enable1(wRegEnTop_6_0), .In1(wRegInTop_6_0), .Enable2(wRegEnBot_6_0), .In2(wRegInBot_6_0), .ScanIn(ScanLink64), .ScanOut(ScanLink63), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_1), .Enable1(wRegEnTop_6_1), .In1(wRegInTop_6_1), .Enable2(wRegEnBot_6_1), .In2(wRegInBot_6_1), .ScanIn(ScanLink65), .ScanOut(ScanLink64), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_2), .Enable1(wRegEnTop_6_2), .In1(wRegInTop_6_2), .Enable2(wRegEnBot_6_2), .In2(wRegInBot_6_2), .ScanIn(ScanLink66), .ScanOut(ScanLink65), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_3), .Enable1(wRegEnTop_6_3), .In1(wRegInTop_6_3), .Enable2(wRegEnBot_6_3), .In2(wRegInBot_6_3), .ScanIn(ScanLink67), .ScanOut(ScanLink66), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_4), .Enable1(wRegEnTop_6_4), .In1(wRegInTop_6_4), .Enable2(wRegEnBot_6_4), .In2(wRegInBot_6_4), .ScanIn(ScanLink68), .ScanOut(ScanLink67), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_5), .Enable1(wRegEnTop_6_5), .In1(wRegInTop_6_5), .Enable2(wRegEnBot_6_5), .In2(wRegInBot_6_5), .ScanIn(ScanLink69), .ScanOut(ScanLink68), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_6), .Enable1(wRegEnTop_6_6), .In1(wRegInTop_6_6), .Enable2(wRegEnBot_6_6), .In2(wRegInBot_6_6), .ScanIn(ScanLink70), .ScanOut(ScanLink69), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_7), .Enable1(wRegEnTop_6_7), .In1(wRegInTop_6_7), .Enable2(wRegEnBot_6_7), .In2(wRegInBot_6_7), .ScanIn(ScanLink71), .ScanOut(ScanLink70), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_8), .Enable1(wRegEnTop_6_8), .In1(wRegInTop_6_8), .Enable2(wRegEnBot_6_8), .In2(wRegInBot_6_8), .ScanIn(ScanLink72), .ScanOut(ScanLink71), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_9), .Enable1(wRegEnTop_6_9), .In1(wRegInTop_6_9), .Enable2(wRegEnBot_6_9), .In2(wRegInBot_6_9), .ScanIn(ScanLink73), .ScanOut(ScanLink72), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_10), .Enable1(wRegEnTop_6_10), .In1(wRegInTop_6_10), .Enable2(wRegEnBot_6_10), .In2(wRegInBot_6_10), .ScanIn(ScanLink74), .ScanOut(ScanLink73), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_11), .Enable1(wRegEnTop_6_11), .In1(wRegInTop_6_11), .Enable2(wRegEnBot_6_11), .In2(wRegInBot_6_11), .ScanIn(ScanLink75), .ScanOut(ScanLink74), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_12), .Enable1(wRegEnTop_6_12), .In1(wRegInTop_6_12), .Enable2(wRegEnBot_6_12), .In2(wRegInBot_6_12), .ScanIn(ScanLink76), .ScanOut(ScanLink75), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_13), .Enable1(wRegEnTop_6_13), .In1(wRegInTop_6_13), .Enable2(wRegEnBot_6_13), .In2(wRegInBot_6_13), .ScanIn(ScanLink77), .ScanOut(ScanLink76), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_14), .Enable1(wRegEnTop_6_14), .In1(wRegInTop_6_14), .Enable2(wRegEnBot_6_14), .In2(wRegInBot_6_14), .ScanIn(ScanLink78), .ScanOut(ScanLink77), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_15), .Enable1(wRegEnTop_6_15), .In1(wRegInTop_6_15), .Enable2(wRegEnBot_6_15), .In2(wRegInBot_6_15), .ScanIn(ScanLink79), .ScanOut(ScanLink78), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_16), .Enable1(wRegEnTop_6_16), .In1(wRegInTop_6_16), .Enable2(wRegEnBot_6_16), .In2(wRegInBot_6_16), .ScanIn(ScanLink80), .ScanOut(ScanLink79), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_17), .Enable1(wRegEnTop_6_17), .In1(wRegInTop_6_17), .Enable2(wRegEnBot_6_17), .In2(wRegInBot_6_17), .ScanIn(ScanLink81), .ScanOut(ScanLink80), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_18), .Enable1(wRegEnTop_6_18), .In1(wRegInTop_6_18), .Enable2(wRegEnBot_6_18), .In2(wRegInBot_6_18), .ScanIn(ScanLink82), .ScanOut(ScanLink81), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_19), .Enable1(wRegEnTop_6_19), .In1(wRegInTop_6_19), .Enable2(wRegEnBot_6_19), .In2(wRegInBot_6_19), .ScanIn(ScanLink83), .ScanOut(ScanLink82), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_20), .Enable1(wRegEnTop_6_20), .In1(wRegInTop_6_20), .Enable2(wRegEnBot_6_20), .In2(wRegInBot_6_20), .ScanIn(ScanLink84), .ScanOut(ScanLink83), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_21), .Enable1(wRegEnTop_6_21), .In1(wRegInTop_6_21), .Enable2(wRegEnBot_6_21), .In2(wRegInBot_6_21), .ScanIn(ScanLink85), .ScanOut(ScanLink84), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_22), .Enable1(wRegEnTop_6_22), .In1(wRegInTop_6_22), .Enable2(wRegEnBot_6_22), .In2(wRegInBot_6_22), .ScanIn(ScanLink86), .ScanOut(ScanLink85), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_23), .Enable1(wRegEnTop_6_23), .In1(wRegInTop_6_23), .Enable2(wRegEnBot_6_23), .In2(wRegInBot_6_23), .ScanIn(ScanLink87), .ScanOut(ScanLink86), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_24), .Enable1(wRegEnTop_6_24), .In1(wRegInTop_6_24), .Enable2(wRegEnBot_6_24), .In2(wRegInBot_6_24), .ScanIn(ScanLink88), .ScanOut(ScanLink87), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_25), .Enable1(wRegEnTop_6_25), .In1(wRegInTop_6_25), .Enable2(wRegEnBot_6_25), .In2(wRegInBot_6_25), .ScanIn(ScanLink89), .ScanOut(ScanLink88), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_26), .Enable1(wRegEnTop_6_26), .In1(wRegInTop_6_26), .Enable2(wRegEnBot_6_26), .In2(wRegInBot_6_26), .ScanIn(ScanLink90), .ScanOut(ScanLink89), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_27), .Enable1(wRegEnTop_6_27), .In1(wRegInTop_6_27), .Enable2(wRegEnBot_6_27), .In2(wRegInBot_6_27), .ScanIn(ScanLink91), .ScanOut(ScanLink90), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_28), .Enable1(wRegEnTop_6_28), .In1(wRegInTop_6_28), .Enable2(wRegEnBot_6_28), .In2(wRegInBot_6_28), .ScanIn(ScanLink92), .ScanOut(ScanLink91), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_29), .Enable1(wRegEnTop_6_29), .In1(wRegInTop_6_29), .Enable2(wRegEnBot_6_29), .In2(wRegInBot_6_29), .ScanIn(ScanLink93), .ScanOut(ScanLink92), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_30), .Enable1(wRegEnTop_6_30), .In1(wRegInTop_6_30), .Enable2(wRegEnBot_6_30), .In2(wRegInBot_6_30), .ScanIn(ScanLink94), .ScanOut(ScanLink93), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_31), .Enable1(wRegEnTop_6_31), .In1(wRegInTop_6_31), .Enable2(wRegEnBot_6_31), .In2(wRegInBot_6_31), .ScanIn(ScanLink95), .ScanOut(ScanLink94), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_32), .Enable1(wRegEnTop_6_32), .In1(wRegInTop_6_32), .Enable2(wRegEnBot_6_32), .In2(wRegInBot_6_32), .ScanIn(ScanLink96), .ScanOut(ScanLink95), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_33), .Enable1(wRegEnTop_6_33), .In1(wRegInTop_6_33), .Enable2(wRegEnBot_6_33), .In2(wRegInBot_6_33), .ScanIn(ScanLink97), .ScanOut(ScanLink96), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_34), .Enable1(wRegEnTop_6_34), .In1(wRegInTop_6_34), .Enable2(wRegEnBot_6_34), .In2(wRegInBot_6_34), .ScanIn(ScanLink98), .ScanOut(ScanLink97), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_35), .Enable1(wRegEnTop_6_35), .In1(wRegInTop_6_35), .Enable2(wRegEnBot_6_35), .In2(wRegInBot_6_35), .ScanIn(ScanLink99), .ScanOut(ScanLink98), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_36), .Enable1(wRegEnTop_6_36), .In1(wRegInTop_6_36), .Enable2(wRegEnBot_6_36), .In2(wRegInBot_6_36), .ScanIn(ScanLink100), .ScanOut(ScanLink99), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_37), .Enable1(wRegEnTop_6_37), .In1(wRegInTop_6_37), .Enable2(wRegEnBot_6_37), .In2(wRegInBot_6_37), .ScanIn(ScanLink101), .ScanOut(ScanLink100), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_38), .Enable1(wRegEnTop_6_38), .In1(wRegInTop_6_38), .Enable2(wRegEnBot_6_38), .In2(wRegInBot_6_38), .ScanIn(ScanLink102), .ScanOut(ScanLink101), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_39), .Enable1(wRegEnTop_6_39), .In1(wRegInTop_6_39), .Enable2(wRegEnBot_6_39), .In2(wRegInBot_6_39), .ScanIn(ScanLink103), .ScanOut(ScanLink102), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_40), .Enable1(wRegEnTop_6_40), .In1(wRegInTop_6_40), .Enable2(wRegEnBot_6_40), .In2(wRegInBot_6_40), .ScanIn(ScanLink104), .ScanOut(ScanLink103), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_41), .Enable1(wRegEnTop_6_41), .In1(wRegInTop_6_41), .Enable2(wRegEnBot_6_41), .In2(wRegInBot_6_41), .ScanIn(ScanLink105), .ScanOut(ScanLink104), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_42), .Enable1(wRegEnTop_6_42), .In1(wRegInTop_6_42), .Enable2(wRegEnBot_6_42), .In2(wRegInBot_6_42), .ScanIn(ScanLink106), .ScanOut(ScanLink105), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_43), .Enable1(wRegEnTop_6_43), .In1(wRegInTop_6_43), .Enable2(wRegEnBot_6_43), .In2(wRegInBot_6_43), .ScanIn(ScanLink107), .ScanOut(ScanLink106), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_44), .Enable1(wRegEnTop_6_44), .In1(wRegInTop_6_44), .Enable2(wRegEnBot_6_44), .In2(wRegInBot_6_44), .ScanIn(ScanLink108), .ScanOut(ScanLink107), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_45), .Enable1(wRegEnTop_6_45), .In1(wRegInTop_6_45), .Enable2(wRegEnBot_6_45), .In2(wRegInBot_6_45), .ScanIn(ScanLink109), .ScanOut(ScanLink108), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_46), .Enable1(wRegEnTop_6_46), .In1(wRegInTop_6_46), .Enable2(wRegEnBot_6_46), .In2(wRegInBot_6_46), .ScanIn(ScanLink110), .ScanOut(ScanLink109), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_47), .Enable1(wRegEnTop_6_47), .In1(wRegInTop_6_47), .Enable2(wRegEnBot_6_47), .In2(wRegInBot_6_47), .ScanIn(ScanLink111), .ScanOut(ScanLink110), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_48), .Enable1(wRegEnTop_6_48), .In1(wRegInTop_6_48), .Enable2(wRegEnBot_6_48), .In2(wRegInBot_6_48), .ScanIn(ScanLink112), .ScanOut(ScanLink111), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_49), .Enable1(wRegEnTop_6_49), .In1(wRegInTop_6_49), .Enable2(wRegEnBot_6_49), .In2(wRegInBot_6_49), .ScanIn(ScanLink113), .ScanOut(ScanLink112), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_50), .Enable1(wRegEnTop_6_50), .In1(wRegInTop_6_50), .Enable2(wRegEnBot_6_50), .In2(wRegInBot_6_50), .ScanIn(ScanLink114), .ScanOut(ScanLink113), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_51), .Enable1(wRegEnTop_6_51), .In1(wRegInTop_6_51), .Enable2(wRegEnBot_6_51), .In2(wRegInBot_6_51), .ScanIn(ScanLink115), .ScanOut(ScanLink114), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_52), .Enable1(wRegEnTop_6_52), .In1(wRegInTop_6_52), .Enable2(wRegEnBot_6_52), .In2(wRegInBot_6_52), .ScanIn(ScanLink116), .ScanOut(ScanLink115), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_53), .Enable1(wRegEnTop_6_53), .In1(wRegInTop_6_53), .Enable2(wRegEnBot_6_53), .In2(wRegInBot_6_53), .ScanIn(ScanLink117), .ScanOut(ScanLink116), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_54), .Enable1(wRegEnTop_6_54), .In1(wRegInTop_6_54), .Enable2(wRegEnBot_6_54), .In2(wRegInBot_6_54), .ScanIn(ScanLink118), .ScanOut(ScanLink117), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_55), .Enable1(wRegEnTop_6_55), .In1(wRegInTop_6_55), .Enable2(wRegEnBot_6_55), .In2(wRegInBot_6_55), .ScanIn(ScanLink119), .ScanOut(ScanLink118), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_56), .Enable1(wRegEnTop_6_56), .In1(wRegInTop_6_56), .Enable2(wRegEnBot_6_56), .In2(wRegInBot_6_56), .ScanIn(ScanLink120), .ScanOut(ScanLink119), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_57), .Enable1(wRegEnTop_6_57), .In1(wRegInTop_6_57), .Enable2(wRegEnBot_6_57), .In2(wRegInBot_6_57), .ScanIn(ScanLink121), .ScanOut(ScanLink120), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_58), .Enable1(wRegEnTop_6_58), .In1(wRegInTop_6_58), .Enable2(wRegEnBot_6_58), .In2(wRegInBot_6_58), .ScanIn(ScanLink122), .ScanOut(ScanLink121), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_59), .Enable1(wRegEnTop_6_59), .In1(wRegInTop_6_59), .Enable2(wRegEnBot_6_59), .In2(wRegInBot_6_59), .ScanIn(ScanLink123), .ScanOut(ScanLink122), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_60), .Enable1(wRegEnTop_6_60), .In1(wRegInTop_6_60), .Enable2(wRegEnBot_6_60), .In2(wRegInBot_6_60), .ScanIn(ScanLink124), .ScanOut(ScanLink123), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_61), .Enable1(wRegEnTop_6_61), .In1(wRegInTop_6_61), .Enable2(wRegEnBot_6_61), .In2(wRegInBot_6_61), .ScanIn(ScanLink125), .ScanOut(ScanLink124), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_62), .Enable1(wRegEnTop_6_62), .In1(wRegInTop_6_62), .Enable2(wRegEnBot_6_62), .In2(wRegInBot_6_62), .ScanIn(ScanLink126), .ScanOut(ScanLink125), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_6_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_6_63), .Enable1(wRegEnTop_6_63), .In1(wRegInTop_6_63), .Enable2(wRegEnBot_6_63), .In2(wRegInBot_6_63), .ScanIn(ScanLink127), .ScanOut(ScanLink126), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_0), .Enable1(wRegEnTop_7_0), .In1(wRegInTop_7_0), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink128), .ScanOut(ScanLink127), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_1), .Enable1(wRegEnTop_7_1), .In1(wRegInTop_7_1), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink129), .ScanOut(ScanLink128), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_2), .Enable1(wRegEnTop_7_2), .In1(wRegInTop_7_2), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink130), .ScanOut(ScanLink129), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_3), .Enable1(wRegEnTop_7_3), .In1(wRegInTop_7_3), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink131), .ScanOut(ScanLink130), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_4), .Enable1(wRegEnTop_7_4), .In1(wRegInTop_7_4), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink132), .ScanOut(ScanLink131), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_5), .Enable1(wRegEnTop_7_5), .In1(wRegInTop_7_5), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink133), .ScanOut(ScanLink132), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_6), .Enable1(wRegEnTop_7_6), .In1(wRegInTop_7_6), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink134), .ScanOut(ScanLink133), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_7), .Enable1(wRegEnTop_7_7), .In1(wRegInTop_7_7), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink135), .ScanOut(ScanLink134), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_8), .Enable1(wRegEnTop_7_8), .In1(wRegInTop_7_8), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink136), .ScanOut(ScanLink135), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_9), .Enable1(wRegEnTop_7_9), .In1(wRegInTop_7_9), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink137), .ScanOut(ScanLink136), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_10), .Enable1(wRegEnTop_7_10), .In1(wRegInTop_7_10), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink138), .ScanOut(ScanLink137), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_11), .Enable1(wRegEnTop_7_11), .In1(wRegInTop_7_11), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink139), .ScanOut(ScanLink138), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_12), .Enable1(wRegEnTop_7_12), .In1(wRegInTop_7_12), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink140), .ScanOut(ScanLink139), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_13), .Enable1(wRegEnTop_7_13), .In1(wRegInTop_7_13), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink141), .ScanOut(ScanLink140), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_14), .Enable1(wRegEnTop_7_14), .In1(wRegInTop_7_14), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink142), .ScanOut(ScanLink141), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_15), .Enable1(wRegEnTop_7_15), .In1(wRegInTop_7_15), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink143), .ScanOut(ScanLink142), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_16), .Enable1(wRegEnTop_7_16), .In1(wRegInTop_7_16), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink144), .ScanOut(ScanLink143), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_17), .Enable1(wRegEnTop_7_17), .In1(wRegInTop_7_17), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink145), .ScanOut(ScanLink144), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_18), .Enable1(wRegEnTop_7_18), .In1(wRegInTop_7_18), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink146), .ScanOut(ScanLink145), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_19), .Enable1(wRegEnTop_7_19), .In1(wRegInTop_7_19), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink147), .ScanOut(ScanLink146), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_20), .Enable1(wRegEnTop_7_20), .In1(wRegInTop_7_20), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink148), .ScanOut(ScanLink147), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_21), .Enable1(wRegEnTop_7_21), .In1(wRegInTop_7_21), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink149), .ScanOut(ScanLink148), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_22), .Enable1(wRegEnTop_7_22), .In1(wRegInTop_7_22), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink150), .ScanOut(ScanLink149), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_23), .Enable1(wRegEnTop_7_23), .In1(wRegInTop_7_23), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink151), .ScanOut(ScanLink150), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_24), .Enable1(wRegEnTop_7_24), .In1(wRegInTop_7_24), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink152), .ScanOut(ScanLink151), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_25), .Enable1(wRegEnTop_7_25), .In1(wRegInTop_7_25), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink153), .ScanOut(ScanLink152), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_26), .Enable1(wRegEnTop_7_26), .In1(wRegInTop_7_26), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink154), .ScanOut(ScanLink153), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_27), .Enable1(wRegEnTop_7_27), .In1(wRegInTop_7_27), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink155), .ScanOut(ScanLink154), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_28), .Enable1(wRegEnTop_7_28), .In1(wRegInTop_7_28), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink156), .ScanOut(ScanLink155), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_29), .Enable1(wRegEnTop_7_29), .In1(wRegInTop_7_29), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink157), .ScanOut(ScanLink156), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_30), .Enable1(wRegEnTop_7_30), .In1(wRegInTop_7_30), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink158), .ScanOut(ScanLink157), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_31), .Enable1(wRegEnTop_7_31), .In1(wRegInTop_7_31), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink159), .ScanOut(ScanLink158), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_32), .Enable1(wRegEnTop_7_32), .In1(wRegInTop_7_32), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink160), .ScanOut(ScanLink159), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_33), .Enable1(wRegEnTop_7_33), .In1(wRegInTop_7_33), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink161), .ScanOut(ScanLink160), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_34), .Enable1(wRegEnTop_7_34), .In1(wRegInTop_7_34), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink162), .ScanOut(ScanLink161), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_35), .Enable1(wRegEnTop_7_35), .In1(wRegInTop_7_35), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink163), .ScanOut(ScanLink162), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_36), .Enable1(wRegEnTop_7_36), .In1(wRegInTop_7_36), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink164), .ScanOut(ScanLink163), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_37), .Enable1(wRegEnTop_7_37), .In1(wRegInTop_7_37), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink165), .ScanOut(ScanLink164), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_38), .Enable1(wRegEnTop_7_38), .In1(wRegInTop_7_38), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink166), .ScanOut(ScanLink165), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_39), .Enable1(wRegEnTop_7_39), .In1(wRegInTop_7_39), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink167), .ScanOut(ScanLink166), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_40), .Enable1(wRegEnTop_7_40), .In1(wRegInTop_7_40), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink168), .ScanOut(ScanLink167), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_41), .Enable1(wRegEnTop_7_41), .In1(wRegInTop_7_41), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink169), .ScanOut(ScanLink168), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_42), .Enable1(wRegEnTop_7_42), .In1(wRegInTop_7_42), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink170), .ScanOut(ScanLink169), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_43), .Enable1(wRegEnTop_7_43), .In1(wRegInTop_7_43), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink171), .ScanOut(ScanLink170), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_44), .Enable1(wRegEnTop_7_44), .In1(wRegInTop_7_44), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink172), .ScanOut(ScanLink171), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_45), .Enable1(wRegEnTop_7_45), .In1(wRegInTop_7_45), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink173), .ScanOut(ScanLink172), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_46), .Enable1(wRegEnTop_7_46), .In1(wRegInTop_7_46), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink174), .ScanOut(ScanLink173), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_47), .Enable1(wRegEnTop_7_47), .In1(wRegInTop_7_47), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink175), .ScanOut(ScanLink174), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_48), .Enable1(wRegEnTop_7_48), .In1(wRegInTop_7_48), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink176), .ScanOut(ScanLink175), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_49), .Enable1(wRegEnTop_7_49), .In1(wRegInTop_7_49), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink177), .ScanOut(ScanLink176), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_50), .Enable1(wRegEnTop_7_50), .In1(wRegInTop_7_50), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink178), .ScanOut(ScanLink177), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_51), .Enable1(wRegEnTop_7_51), .In1(wRegInTop_7_51), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink179), .ScanOut(ScanLink178), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_52), .Enable1(wRegEnTop_7_52), .In1(wRegInTop_7_52), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink180), .ScanOut(ScanLink179), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_53), .Enable1(wRegEnTop_7_53), .In1(wRegInTop_7_53), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink181), .ScanOut(ScanLink180), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_54), .Enable1(wRegEnTop_7_54), .In1(wRegInTop_7_54), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink182), .ScanOut(ScanLink181), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_55), .Enable1(wRegEnTop_7_55), .In1(wRegInTop_7_55), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink183), .ScanOut(ScanLink182), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_56), .Enable1(wRegEnTop_7_56), .In1(wRegInTop_7_56), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink184), .ScanOut(ScanLink183), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_57), .Enable1(wRegEnTop_7_57), .In1(wRegInTop_7_57), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink185), .ScanOut(ScanLink184), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_58), .Enable1(wRegEnTop_7_58), .In1(wRegInTop_7_58), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink186), .ScanOut(ScanLink185), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_59), .Enable1(wRegEnTop_7_59), .In1(wRegInTop_7_59), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink187), .ScanOut(ScanLink186), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_60), .Enable1(wRegEnTop_7_60), .In1(wRegInTop_7_60), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink188), .ScanOut(ScanLink187), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_61), .Enable1(wRegEnTop_7_61), .In1(wRegInTop_7_61), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink189), .ScanOut(ScanLink188), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_62), .Enable1(wRegEnTop_7_62), .In1(wRegInTop_7_62), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink190), .ScanOut(ScanLink189), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_63), .Enable1(wRegEnTop_7_63), .In1(wRegInTop_7_63), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink191), .ScanOut(ScanLink190), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_64), .Enable1(wRegEnTop_7_64), .In1(wRegInTop_7_64), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink192), .ScanOut(ScanLink191), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_65), .Enable1(wRegEnTop_7_65), .In1(wRegInTop_7_65), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink193), .ScanOut(ScanLink192), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_66), .Enable1(wRegEnTop_7_66), .In1(wRegInTop_7_66), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink194), .ScanOut(ScanLink193), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_67), .Enable1(wRegEnTop_7_67), .In1(wRegInTop_7_67), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink195), .ScanOut(ScanLink194), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_68), .Enable1(wRegEnTop_7_68), .In1(wRegInTop_7_68), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink196), .ScanOut(ScanLink195), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_69), .Enable1(wRegEnTop_7_69), .In1(wRegInTop_7_69), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink197), .ScanOut(ScanLink196), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_70), .Enable1(wRegEnTop_7_70), .In1(wRegInTop_7_70), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink198), .ScanOut(ScanLink197), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_71), .Enable1(wRegEnTop_7_71), .In1(wRegInTop_7_71), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink199), .ScanOut(ScanLink198), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_72), .Enable1(wRegEnTop_7_72), .In1(wRegInTop_7_72), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink200), .ScanOut(ScanLink199), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_73), .Enable1(wRegEnTop_7_73), .In1(wRegInTop_7_73), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink201), .ScanOut(ScanLink200), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_74), .Enable1(wRegEnTop_7_74), .In1(wRegInTop_7_74), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink202), .ScanOut(ScanLink201), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_75), .Enable1(wRegEnTop_7_75), .In1(wRegInTop_7_75), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink203), .ScanOut(ScanLink202), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_76), .Enable1(wRegEnTop_7_76), .In1(wRegInTop_7_76), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink204), .ScanOut(ScanLink203), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_77), .Enable1(wRegEnTop_7_77), .In1(wRegInTop_7_77), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink205), .ScanOut(ScanLink204), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_78), .Enable1(wRegEnTop_7_78), .In1(wRegInTop_7_78), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink206), .ScanOut(ScanLink205), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_79), .Enable1(wRegEnTop_7_79), .In1(wRegInTop_7_79), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink207), .ScanOut(ScanLink206), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_80), .Enable1(wRegEnTop_7_80), .In1(wRegInTop_7_80), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink208), .ScanOut(ScanLink207), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_81), .Enable1(wRegEnTop_7_81), .In1(wRegInTop_7_81), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink209), .ScanOut(ScanLink208), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_82), .Enable1(wRegEnTop_7_82), .In1(wRegInTop_7_82), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink210), .ScanOut(ScanLink209), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_83), .Enable1(wRegEnTop_7_83), .In1(wRegInTop_7_83), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink211), .ScanOut(ScanLink210), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_84), .Enable1(wRegEnTop_7_84), .In1(wRegInTop_7_84), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink212), .ScanOut(ScanLink211), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_85), .Enable1(wRegEnTop_7_85), .In1(wRegInTop_7_85), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink213), .ScanOut(ScanLink212), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_86), .Enable1(wRegEnTop_7_86), .In1(wRegInTop_7_86), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink214), .ScanOut(ScanLink213), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_87), .Enable1(wRegEnTop_7_87), .In1(wRegInTop_7_87), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink215), .ScanOut(ScanLink214), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_88), .Enable1(wRegEnTop_7_88), .In1(wRegInTop_7_88), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink216), .ScanOut(ScanLink215), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_89), .Enable1(wRegEnTop_7_89), .In1(wRegInTop_7_89), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink217), .ScanOut(ScanLink216), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_90), .Enable1(wRegEnTop_7_90), .In1(wRegInTop_7_90), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink218), .ScanOut(ScanLink217), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_91), .Enable1(wRegEnTop_7_91), .In1(wRegInTop_7_91), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink219), .ScanOut(ScanLink218), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_92), .Enable1(wRegEnTop_7_92), .In1(wRegInTop_7_92), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink220), .ScanOut(ScanLink219), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_93), .Enable1(wRegEnTop_7_93), .In1(wRegInTop_7_93), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink221), .ScanOut(ScanLink220), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_94), .Enable1(wRegEnTop_7_94), .In1(wRegInTop_7_94), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink222), .ScanOut(ScanLink221), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_95), .Enable1(wRegEnTop_7_95), .In1(wRegInTop_7_95), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink223), .ScanOut(ScanLink222), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_96), .Enable1(wRegEnTop_7_96), .In1(wRegInTop_7_96), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink224), .ScanOut(ScanLink223), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_97), .Enable1(wRegEnTop_7_97), .In1(wRegInTop_7_97), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink225), .ScanOut(ScanLink224), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_98), .Enable1(wRegEnTop_7_98), .In1(wRegInTop_7_98), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink226), .ScanOut(ScanLink225), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_99), .Enable1(wRegEnTop_7_99), .In1(wRegInTop_7_99), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink227), .ScanOut(ScanLink226), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_100), .Enable1(wRegEnTop_7_100), .In1(wRegInTop_7_100), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink228), .ScanOut(ScanLink227), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_101), .Enable1(wRegEnTop_7_101), .In1(wRegInTop_7_101), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink229), .ScanOut(ScanLink228), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_102), .Enable1(wRegEnTop_7_102), .In1(wRegInTop_7_102), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink230), .ScanOut(ScanLink229), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_103), .Enable1(wRegEnTop_7_103), .In1(wRegInTop_7_103), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink231), .ScanOut(ScanLink230), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_104), .Enable1(wRegEnTop_7_104), .In1(wRegInTop_7_104), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink232), .ScanOut(ScanLink231), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_105), .Enable1(wRegEnTop_7_105), .In1(wRegInTop_7_105), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink233), .ScanOut(ScanLink232), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_106), .Enable1(wRegEnTop_7_106), .In1(wRegInTop_7_106), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink234), .ScanOut(ScanLink233), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_107), .Enable1(wRegEnTop_7_107), .In1(wRegInTop_7_107), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink235), .ScanOut(ScanLink234), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_108), .Enable1(wRegEnTop_7_108), .In1(wRegInTop_7_108), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink236), .ScanOut(ScanLink235), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_109), .Enable1(wRegEnTop_7_109), .In1(wRegInTop_7_109), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink237), .ScanOut(ScanLink236), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_110), .Enable1(wRegEnTop_7_110), .In1(wRegInTop_7_110), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink238), .ScanOut(ScanLink237), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_111), .Enable1(wRegEnTop_7_111), .In1(wRegInTop_7_111), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink239), .ScanOut(ScanLink238), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_112), .Enable1(wRegEnTop_7_112), .In1(wRegInTop_7_112), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink240), .ScanOut(ScanLink239), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_113), .Enable1(wRegEnTop_7_113), .In1(wRegInTop_7_113), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink241), .ScanOut(ScanLink240), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_114), .Enable1(wRegEnTop_7_114), .In1(wRegInTop_7_114), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink242), .ScanOut(ScanLink241), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_115), .Enable1(wRegEnTop_7_115), .In1(wRegInTop_7_115), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink243), .ScanOut(ScanLink242), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_116), .Enable1(wRegEnTop_7_116), .In1(wRegInTop_7_116), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink244), .ScanOut(ScanLink243), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_117), .Enable1(wRegEnTop_7_117), .In1(wRegInTop_7_117), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink245), .ScanOut(ScanLink244), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_118), .Enable1(wRegEnTop_7_118), .In1(wRegInTop_7_118), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink246), .ScanOut(ScanLink245), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_119), .Enable1(wRegEnTop_7_119), .In1(wRegInTop_7_119), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink247), .ScanOut(ScanLink246), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_120), .Enable1(wRegEnTop_7_120), .In1(wRegInTop_7_120), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink248), .ScanOut(ScanLink247), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_121), .Enable1(wRegEnTop_7_121), .In1(wRegInTop_7_121), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink249), .ScanOut(ScanLink248), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_122), .Enable1(wRegEnTop_7_122), .In1(wRegInTop_7_122), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink250), .ScanOut(ScanLink249), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_123), .Enable1(wRegEnTop_7_123), .In1(wRegInTop_7_123), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink251), .ScanOut(ScanLink250), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_124), .Enable1(wRegEnTop_7_124), .In1(wRegInTop_7_124), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink252), .ScanOut(ScanLink251), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_125), .Enable1(wRegEnTop_7_125), .In1(wRegInTop_7_125), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink253), .ScanOut(ScanLink252), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_126), .Enable1(wRegEnTop_7_126), .In1(wRegInTop_7_126), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink254), .ScanOut(ScanLink253), .ScanEnable(ScanEnable) );
BHeap_Reg #( 32, 1, 1 ) BHR_7_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(wRegOut_7_127), .Enable1(wRegEnTop_7_127), .In1(wRegInTop_7_127), .Enable2(1'b0), .In2(32'b0), .ScanIn(ScanLink255), .ScanOut(ScanLink254), .ScanEnable(ScanEnable) );
BHeap_Node #( 32 ) BHN_0_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_0), .P_WR(wRegEnBot_0_0), .P_In(wRegOut_0_0), .P_Out(wRegInBot_0_0), .L_WR(wRegEnTop_1_0), .L_In(wRegOut_1_0), .L_Out(wRegInTop_1_0), .R_WR(wRegEnTop_1_1), .R_In(wRegOut_1_1), .R_Out(wRegInTop_1_1) );
BHeap_Node #( 32 ) BHN_1_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_1), .P_WR(wRegEnBot_1_0), .P_In(wRegOut_1_0), .P_Out(wRegInBot_1_0), .L_WR(wRegEnTop_2_0), .L_In(wRegOut_2_0), .L_Out(wRegInTop_2_0), .R_WR(wRegEnTop_2_1), .R_In(wRegOut_2_1), .R_Out(wRegInTop_2_1) );
BHeap_Node #( 32 ) BHN_1_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_1), .P_WR(wRegEnBot_1_1), .P_In(wRegOut_1_1), .P_Out(wRegInBot_1_1), .L_WR(wRegEnTop_2_2), .L_In(wRegOut_2_2), .L_Out(wRegInTop_2_2), .R_WR(wRegEnTop_2_3), .R_In(wRegOut_2_3), .R_Out(wRegInTop_2_3) );
BHeap_Node #( 32 ) BHN_2_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_2), .P_WR(wRegEnBot_2_0), .P_In(wRegOut_2_0), .P_Out(wRegInBot_2_0), .L_WR(wRegEnTop_3_0), .L_In(wRegOut_3_0), .L_Out(wRegInTop_3_0), .R_WR(wRegEnTop_3_1), .R_In(wRegOut_3_1), .R_Out(wRegInTop_3_1) );
BHeap_Node #( 32 ) BHN_2_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_2), .P_WR(wRegEnBot_2_1), .P_In(wRegOut_2_1), .P_Out(wRegInBot_2_1), .L_WR(wRegEnTop_3_2), .L_In(wRegOut_3_2), .L_Out(wRegInTop_3_2), .R_WR(wRegEnTop_3_3), .R_In(wRegOut_3_3), .R_Out(wRegInTop_3_3) );
BHeap_Node #( 32 ) BHN_2_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_2), .P_WR(wRegEnBot_2_2), .P_In(wRegOut_2_2), .P_Out(wRegInBot_2_2), .L_WR(wRegEnTop_3_4), .L_In(wRegOut_3_4), .L_Out(wRegInTop_3_4), .R_WR(wRegEnTop_3_5), .R_In(wRegOut_3_5), .R_Out(wRegInTop_3_5) );
BHeap_Node #( 32 ) BHN_2_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_2), .P_WR(wRegEnBot_2_3), .P_In(wRegOut_2_3), .P_Out(wRegInBot_2_3), .L_WR(wRegEnTop_3_6), .L_In(wRegOut_3_6), .L_Out(wRegInTop_3_6), .R_WR(wRegEnTop_3_7), .R_In(wRegOut_3_7), .R_Out(wRegInTop_3_7) );
BHeap_Node #( 32 ) BHN_3_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_0), .P_In(wRegOut_3_0), .P_Out(wRegInBot_3_0), .L_WR(wRegEnTop_4_0), .L_In(wRegOut_4_0), .L_Out(wRegInTop_4_0), .R_WR(wRegEnTop_4_1), .R_In(wRegOut_4_1), .R_Out(wRegInTop_4_1) );
BHeap_Node #( 32 ) BHN_3_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_1), .P_In(wRegOut_3_1), .P_Out(wRegInBot_3_1), .L_WR(wRegEnTop_4_2), .L_In(wRegOut_4_2), .L_Out(wRegInTop_4_2), .R_WR(wRegEnTop_4_3), .R_In(wRegOut_4_3), .R_Out(wRegInTop_4_3) );
BHeap_Node #( 32 ) BHN_3_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_2), .P_In(wRegOut_3_2), .P_Out(wRegInBot_3_2), .L_WR(wRegEnTop_4_4), .L_In(wRegOut_4_4), .L_Out(wRegInTop_4_4), .R_WR(wRegEnTop_4_5), .R_In(wRegOut_4_5), .R_Out(wRegInTop_4_5) );
BHeap_Node #( 32 ) BHN_3_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_3), .P_In(wRegOut_3_3), .P_Out(wRegInBot_3_3), .L_WR(wRegEnTop_4_6), .L_In(wRegOut_4_6), .L_Out(wRegInTop_4_6), .R_WR(wRegEnTop_4_7), .R_In(wRegOut_4_7), .R_Out(wRegInTop_4_7) );
BHeap_Node #( 32 ) BHN_3_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_4), .P_In(wRegOut_3_4), .P_Out(wRegInBot_3_4), .L_WR(wRegEnTop_4_8), .L_In(wRegOut_4_8), .L_Out(wRegInTop_4_8), .R_WR(wRegEnTop_4_9), .R_In(wRegOut_4_9), .R_Out(wRegInTop_4_9) );
BHeap_Node #( 32 ) BHN_3_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_5), .P_In(wRegOut_3_5), .P_Out(wRegInBot_3_5), .L_WR(wRegEnTop_4_10), .L_In(wRegOut_4_10), .L_Out(wRegInTop_4_10), .R_WR(wRegEnTop_4_11), .R_In(wRegOut_4_11), .R_Out(wRegInTop_4_11) );
BHeap_Node #( 32 ) BHN_3_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_6), .P_In(wRegOut_3_6), .P_Out(wRegInBot_3_6), .L_WR(wRegEnTop_4_12), .L_In(wRegOut_4_12), .L_Out(wRegInTop_4_12), .R_WR(wRegEnTop_4_13), .R_In(wRegOut_4_13), .R_Out(wRegInTop_4_13) );
BHeap_Node #( 32 ) BHN_3_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_3), .P_WR(wRegEnBot_3_7), .P_In(wRegOut_3_7), .P_Out(wRegInBot_3_7), .L_WR(wRegEnTop_4_14), .L_In(wRegOut_4_14), .L_Out(wRegInTop_4_14), .R_WR(wRegEnTop_4_15), .R_In(wRegOut_4_15), .R_Out(wRegInTop_4_15) );
BHeap_Node #( 32 ) BHN_4_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_0), .P_In(wRegOut_4_0), .P_Out(wRegInBot_4_0), .L_WR(wRegEnTop_5_0), .L_In(wRegOut_5_0), .L_Out(wRegInTop_5_0), .R_WR(wRegEnTop_5_1), .R_In(wRegOut_5_1), .R_Out(wRegInTop_5_1) );
BHeap_Node #( 32 ) BHN_4_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_1), .P_In(wRegOut_4_1), .P_Out(wRegInBot_4_1), .L_WR(wRegEnTop_5_2), .L_In(wRegOut_5_2), .L_Out(wRegInTop_5_2), .R_WR(wRegEnTop_5_3), .R_In(wRegOut_5_3), .R_Out(wRegInTop_5_3) );
BHeap_Node #( 32 ) BHN_4_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_2), .P_In(wRegOut_4_2), .P_Out(wRegInBot_4_2), .L_WR(wRegEnTop_5_4), .L_In(wRegOut_5_4), .L_Out(wRegInTop_5_4), .R_WR(wRegEnTop_5_5), .R_In(wRegOut_5_5), .R_Out(wRegInTop_5_5) );
BHeap_Node #( 32 ) BHN_4_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_3), .P_In(wRegOut_4_3), .P_Out(wRegInBot_4_3), .L_WR(wRegEnTop_5_6), .L_In(wRegOut_5_6), .L_Out(wRegInTop_5_6), .R_WR(wRegEnTop_5_7), .R_In(wRegOut_5_7), .R_Out(wRegInTop_5_7) );
BHeap_Node #( 32 ) BHN_4_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_4), .P_In(wRegOut_4_4), .P_Out(wRegInBot_4_4), .L_WR(wRegEnTop_5_8), .L_In(wRegOut_5_8), .L_Out(wRegInTop_5_8), .R_WR(wRegEnTop_5_9), .R_In(wRegOut_5_9), .R_Out(wRegInTop_5_9) );
BHeap_Node #( 32 ) BHN_4_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_5), .P_In(wRegOut_4_5), .P_Out(wRegInBot_4_5), .L_WR(wRegEnTop_5_10), .L_In(wRegOut_5_10), .L_Out(wRegInTop_5_10), .R_WR(wRegEnTop_5_11), .R_In(wRegOut_5_11), .R_Out(wRegInTop_5_11) );
BHeap_Node #( 32 ) BHN_4_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_6), .P_In(wRegOut_4_6), .P_Out(wRegInBot_4_6), .L_WR(wRegEnTop_5_12), .L_In(wRegOut_5_12), .L_Out(wRegInTop_5_12), .R_WR(wRegEnTop_5_13), .R_In(wRegOut_5_13), .R_Out(wRegInTop_5_13) );
BHeap_Node #( 32 ) BHN_4_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_7), .P_In(wRegOut_4_7), .P_Out(wRegInBot_4_7), .L_WR(wRegEnTop_5_14), .L_In(wRegOut_5_14), .L_Out(wRegInTop_5_14), .R_WR(wRegEnTop_5_15), .R_In(wRegOut_5_15), .R_Out(wRegInTop_5_15) );
BHeap_Node #( 32 ) BHN_4_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_8), .P_In(wRegOut_4_8), .P_Out(wRegInBot_4_8), .L_WR(wRegEnTop_5_16), .L_In(wRegOut_5_16), .L_Out(wRegInTop_5_16), .R_WR(wRegEnTop_5_17), .R_In(wRegOut_5_17), .R_Out(wRegInTop_5_17) );
BHeap_Node #( 32 ) BHN_4_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_9), .P_In(wRegOut_4_9), .P_Out(wRegInBot_4_9), .L_WR(wRegEnTop_5_18), .L_In(wRegOut_5_18), .L_Out(wRegInTop_5_18), .R_WR(wRegEnTop_5_19), .R_In(wRegOut_5_19), .R_Out(wRegInTop_5_19) );
BHeap_Node #( 32 ) BHN_4_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_10), .P_In(wRegOut_4_10), .P_Out(wRegInBot_4_10), .L_WR(wRegEnTop_5_20), .L_In(wRegOut_5_20), .L_Out(wRegInTop_5_20), .R_WR(wRegEnTop_5_21), .R_In(wRegOut_5_21), .R_Out(wRegInTop_5_21) );
BHeap_Node #( 32 ) BHN_4_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_11), .P_In(wRegOut_4_11), .P_Out(wRegInBot_4_11), .L_WR(wRegEnTop_5_22), .L_In(wRegOut_5_22), .L_Out(wRegInTop_5_22), .R_WR(wRegEnTop_5_23), .R_In(wRegOut_5_23), .R_Out(wRegInTop_5_23) );
BHeap_Node #( 32 ) BHN_4_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_12), .P_In(wRegOut_4_12), .P_Out(wRegInBot_4_12), .L_WR(wRegEnTop_5_24), .L_In(wRegOut_5_24), .L_Out(wRegInTop_5_24), .R_WR(wRegEnTop_5_25), .R_In(wRegOut_5_25), .R_Out(wRegInTop_5_25) );
BHeap_Node #( 32 ) BHN_4_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_13), .P_In(wRegOut_4_13), .P_Out(wRegInBot_4_13), .L_WR(wRegEnTop_5_26), .L_In(wRegOut_5_26), .L_Out(wRegInTop_5_26), .R_WR(wRegEnTop_5_27), .R_In(wRegOut_5_27), .R_Out(wRegInTop_5_27) );
BHeap_Node #( 32 ) BHN_4_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_14), .P_In(wRegOut_4_14), .P_Out(wRegInBot_4_14), .L_WR(wRegEnTop_5_28), .L_In(wRegOut_5_28), .L_Out(wRegInTop_5_28), .R_WR(wRegEnTop_5_29), .R_In(wRegOut_5_29), .R_Out(wRegInTop_5_29) );
BHeap_Node #( 32 ) BHN_4_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_4), .P_WR(wRegEnBot_4_15), .P_In(wRegOut_4_15), .P_Out(wRegInBot_4_15), .L_WR(wRegEnTop_5_30), .L_In(wRegOut_5_30), .L_Out(wRegInTop_5_30), .R_WR(wRegEnTop_5_31), .R_In(wRegOut_5_31), .R_Out(wRegInTop_5_31) );
BHeap_Node #( 32 ) BHN_5_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_0), .P_In(wRegOut_5_0), .P_Out(wRegInBot_5_0), .L_WR(wRegEnTop_6_0), .L_In(wRegOut_6_0), .L_Out(wRegInTop_6_0), .R_WR(wRegEnTop_6_1), .R_In(wRegOut_6_1), .R_Out(wRegInTop_6_1) );
BHeap_Node #( 32 ) BHN_5_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_1), .P_In(wRegOut_5_1), .P_Out(wRegInBot_5_1), .L_WR(wRegEnTop_6_2), .L_In(wRegOut_6_2), .L_Out(wRegInTop_6_2), .R_WR(wRegEnTop_6_3), .R_In(wRegOut_6_3), .R_Out(wRegInTop_6_3) );
BHeap_Node #( 32 ) BHN_5_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_2), .P_In(wRegOut_5_2), .P_Out(wRegInBot_5_2), .L_WR(wRegEnTop_6_4), .L_In(wRegOut_6_4), .L_Out(wRegInTop_6_4), .R_WR(wRegEnTop_6_5), .R_In(wRegOut_6_5), .R_Out(wRegInTop_6_5) );
BHeap_Node #( 32 ) BHN_5_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_3), .P_In(wRegOut_5_3), .P_Out(wRegInBot_5_3), .L_WR(wRegEnTop_6_6), .L_In(wRegOut_6_6), .L_Out(wRegInTop_6_6), .R_WR(wRegEnTop_6_7), .R_In(wRegOut_6_7), .R_Out(wRegInTop_6_7) );
BHeap_Node #( 32 ) BHN_5_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_4), .P_In(wRegOut_5_4), .P_Out(wRegInBot_5_4), .L_WR(wRegEnTop_6_8), .L_In(wRegOut_6_8), .L_Out(wRegInTop_6_8), .R_WR(wRegEnTop_6_9), .R_In(wRegOut_6_9), .R_Out(wRegInTop_6_9) );
BHeap_Node #( 32 ) BHN_5_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_5), .P_In(wRegOut_5_5), .P_Out(wRegInBot_5_5), .L_WR(wRegEnTop_6_10), .L_In(wRegOut_6_10), .L_Out(wRegInTop_6_10), .R_WR(wRegEnTop_6_11), .R_In(wRegOut_6_11), .R_Out(wRegInTop_6_11) );
BHeap_Node #( 32 ) BHN_5_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_6), .P_In(wRegOut_5_6), .P_Out(wRegInBot_5_6), .L_WR(wRegEnTop_6_12), .L_In(wRegOut_6_12), .L_Out(wRegInTop_6_12), .R_WR(wRegEnTop_6_13), .R_In(wRegOut_6_13), .R_Out(wRegInTop_6_13) );
BHeap_Node #( 32 ) BHN_5_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_7), .P_In(wRegOut_5_7), .P_Out(wRegInBot_5_7), .L_WR(wRegEnTop_6_14), .L_In(wRegOut_6_14), .L_Out(wRegInTop_6_14), .R_WR(wRegEnTop_6_15), .R_In(wRegOut_6_15), .R_Out(wRegInTop_6_15) );
BHeap_Node #( 32 ) BHN_5_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_8), .P_In(wRegOut_5_8), .P_Out(wRegInBot_5_8), .L_WR(wRegEnTop_6_16), .L_In(wRegOut_6_16), .L_Out(wRegInTop_6_16), .R_WR(wRegEnTop_6_17), .R_In(wRegOut_6_17), .R_Out(wRegInTop_6_17) );
BHeap_Node #( 32 ) BHN_5_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_9), .P_In(wRegOut_5_9), .P_Out(wRegInBot_5_9), .L_WR(wRegEnTop_6_18), .L_In(wRegOut_6_18), .L_Out(wRegInTop_6_18), .R_WR(wRegEnTop_6_19), .R_In(wRegOut_6_19), .R_Out(wRegInTop_6_19) );
BHeap_Node #( 32 ) BHN_5_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_10), .P_In(wRegOut_5_10), .P_Out(wRegInBot_5_10), .L_WR(wRegEnTop_6_20), .L_In(wRegOut_6_20), .L_Out(wRegInTop_6_20), .R_WR(wRegEnTop_6_21), .R_In(wRegOut_6_21), .R_Out(wRegInTop_6_21) );
BHeap_Node #( 32 ) BHN_5_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_11), .P_In(wRegOut_5_11), .P_Out(wRegInBot_5_11), .L_WR(wRegEnTop_6_22), .L_In(wRegOut_6_22), .L_Out(wRegInTop_6_22), .R_WR(wRegEnTop_6_23), .R_In(wRegOut_6_23), .R_Out(wRegInTop_6_23) );
BHeap_Node #( 32 ) BHN_5_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_12), .P_In(wRegOut_5_12), .P_Out(wRegInBot_5_12), .L_WR(wRegEnTop_6_24), .L_In(wRegOut_6_24), .L_Out(wRegInTop_6_24), .R_WR(wRegEnTop_6_25), .R_In(wRegOut_6_25), .R_Out(wRegInTop_6_25) );
BHeap_Node #( 32 ) BHN_5_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_13), .P_In(wRegOut_5_13), .P_Out(wRegInBot_5_13), .L_WR(wRegEnTop_6_26), .L_In(wRegOut_6_26), .L_Out(wRegInTop_6_26), .R_WR(wRegEnTop_6_27), .R_In(wRegOut_6_27), .R_Out(wRegInTop_6_27) );
BHeap_Node #( 32 ) BHN_5_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_14), .P_In(wRegOut_5_14), .P_Out(wRegInBot_5_14), .L_WR(wRegEnTop_6_28), .L_In(wRegOut_6_28), .L_Out(wRegInTop_6_28), .R_WR(wRegEnTop_6_29), .R_In(wRegOut_6_29), .R_Out(wRegInTop_6_29) );
BHeap_Node #( 32 ) BHN_5_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_15), .P_In(wRegOut_5_15), .P_Out(wRegInBot_5_15), .L_WR(wRegEnTop_6_30), .L_In(wRegOut_6_30), .L_Out(wRegInTop_6_30), .R_WR(wRegEnTop_6_31), .R_In(wRegOut_6_31), .R_Out(wRegInTop_6_31) );
BHeap_Node #( 32 ) BHN_5_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_16), .P_In(wRegOut_5_16), .P_Out(wRegInBot_5_16), .L_WR(wRegEnTop_6_32), .L_In(wRegOut_6_32), .L_Out(wRegInTop_6_32), .R_WR(wRegEnTop_6_33), .R_In(wRegOut_6_33), .R_Out(wRegInTop_6_33) );
BHeap_Node #( 32 ) BHN_5_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_17), .P_In(wRegOut_5_17), .P_Out(wRegInBot_5_17), .L_WR(wRegEnTop_6_34), .L_In(wRegOut_6_34), .L_Out(wRegInTop_6_34), .R_WR(wRegEnTop_6_35), .R_In(wRegOut_6_35), .R_Out(wRegInTop_6_35) );
BHeap_Node #( 32 ) BHN_5_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_18), .P_In(wRegOut_5_18), .P_Out(wRegInBot_5_18), .L_WR(wRegEnTop_6_36), .L_In(wRegOut_6_36), .L_Out(wRegInTop_6_36), .R_WR(wRegEnTop_6_37), .R_In(wRegOut_6_37), .R_Out(wRegInTop_6_37) );
BHeap_Node #( 32 ) BHN_5_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_19), .P_In(wRegOut_5_19), .P_Out(wRegInBot_5_19), .L_WR(wRegEnTop_6_38), .L_In(wRegOut_6_38), .L_Out(wRegInTop_6_38), .R_WR(wRegEnTop_6_39), .R_In(wRegOut_6_39), .R_Out(wRegInTop_6_39) );
BHeap_Node #( 32 ) BHN_5_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_20), .P_In(wRegOut_5_20), .P_Out(wRegInBot_5_20), .L_WR(wRegEnTop_6_40), .L_In(wRegOut_6_40), .L_Out(wRegInTop_6_40), .R_WR(wRegEnTop_6_41), .R_In(wRegOut_6_41), .R_Out(wRegInTop_6_41) );
BHeap_Node #( 32 ) BHN_5_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_21), .P_In(wRegOut_5_21), .P_Out(wRegInBot_5_21), .L_WR(wRegEnTop_6_42), .L_In(wRegOut_6_42), .L_Out(wRegInTop_6_42), .R_WR(wRegEnTop_6_43), .R_In(wRegOut_6_43), .R_Out(wRegInTop_6_43) );
BHeap_Node #( 32 ) BHN_5_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_22), .P_In(wRegOut_5_22), .P_Out(wRegInBot_5_22), .L_WR(wRegEnTop_6_44), .L_In(wRegOut_6_44), .L_Out(wRegInTop_6_44), .R_WR(wRegEnTop_6_45), .R_In(wRegOut_6_45), .R_Out(wRegInTop_6_45) );
BHeap_Node #( 32 ) BHN_5_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_23), .P_In(wRegOut_5_23), .P_Out(wRegInBot_5_23), .L_WR(wRegEnTop_6_46), .L_In(wRegOut_6_46), .L_Out(wRegInTop_6_46), .R_WR(wRegEnTop_6_47), .R_In(wRegOut_6_47), .R_Out(wRegInTop_6_47) );
BHeap_Node #( 32 ) BHN_5_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_24), .P_In(wRegOut_5_24), .P_Out(wRegInBot_5_24), .L_WR(wRegEnTop_6_48), .L_In(wRegOut_6_48), .L_Out(wRegInTop_6_48), .R_WR(wRegEnTop_6_49), .R_In(wRegOut_6_49), .R_Out(wRegInTop_6_49) );
BHeap_Node #( 32 ) BHN_5_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_25), .P_In(wRegOut_5_25), .P_Out(wRegInBot_5_25), .L_WR(wRegEnTop_6_50), .L_In(wRegOut_6_50), .L_Out(wRegInTop_6_50), .R_WR(wRegEnTop_6_51), .R_In(wRegOut_6_51), .R_Out(wRegInTop_6_51) );
BHeap_Node #( 32 ) BHN_5_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_26), .P_In(wRegOut_5_26), .P_Out(wRegInBot_5_26), .L_WR(wRegEnTop_6_52), .L_In(wRegOut_6_52), .L_Out(wRegInTop_6_52), .R_WR(wRegEnTop_6_53), .R_In(wRegOut_6_53), .R_Out(wRegInTop_6_53) );
BHeap_Node #( 32 ) BHN_5_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_27), .P_In(wRegOut_5_27), .P_Out(wRegInBot_5_27), .L_WR(wRegEnTop_6_54), .L_In(wRegOut_6_54), .L_Out(wRegInTop_6_54), .R_WR(wRegEnTop_6_55), .R_In(wRegOut_6_55), .R_Out(wRegInTop_6_55) );
BHeap_Node #( 32 ) BHN_5_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_28), .P_In(wRegOut_5_28), .P_Out(wRegInBot_5_28), .L_WR(wRegEnTop_6_56), .L_In(wRegOut_6_56), .L_Out(wRegInTop_6_56), .R_WR(wRegEnTop_6_57), .R_In(wRegOut_6_57), .R_Out(wRegInTop_6_57) );
BHeap_Node #( 32 ) BHN_5_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_29), .P_In(wRegOut_5_29), .P_Out(wRegInBot_5_29), .L_WR(wRegEnTop_6_58), .L_In(wRegOut_6_58), .L_Out(wRegInTop_6_58), .R_WR(wRegEnTop_6_59), .R_In(wRegOut_6_59), .R_Out(wRegInTop_6_59) );
BHeap_Node #( 32 ) BHN_5_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_30), .P_In(wRegOut_5_30), .P_Out(wRegInBot_5_30), .L_WR(wRegEnTop_6_60), .L_In(wRegOut_6_60), .L_Out(wRegInTop_6_60), .R_WR(wRegEnTop_6_61), .R_In(wRegOut_6_61), .R_Out(wRegInTop_6_61) );
BHeap_Node #( 32 ) BHN_5_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_5), .P_WR(wRegEnBot_5_31), .P_In(wRegOut_5_31), .P_Out(wRegInBot_5_31), .L_WR(wRegEnTop_6_62), .L_In(wRegOut_6_62), .L_Out(wRegInTop_6_62), .R_WR(wRegEnTop_6_63), .R_In(wRegOut_6_63), .R_Out(wRegInTop_6_63) );
BHeap_Node #( 32 ) BHN_6_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_0), .P_In(wRegOut_6_0), .P_Out(wRegInBot_6_0), .L_WR(wRegEnTop_7_0), .L_In(wRegOut_7_0), .L_Out(wRegInTop_7_0), .R_WR(wRegEnTop_7_1), .R_In(wRegOut_7_1), .R_Out(wRegInTop_7_1) );
BHeap_Node #( 32 ) BHN_6_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_1), .P_In(wRegOut_6_1), .P_Out(wRegInBot_6_1), .L_WR(wRegEnTop_7_2), .L_In(wRegOut_7_2), .L_Out(wRegInTop_7_2), .R_WR(wRegEnTop_7_3), .R_In(wRegOut_7_3), .R_Out(wRegInTop_7_3) );
BHeap_Node #( 32 ) BHN_6_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_2), .P_In(wRegOut_6_2), .P_Out(wRegInBot_6_2), .L_WR(wRegEnTop_7_4), .L_In(wRegOut_7_4), .L_Out(wRegInTop_7_4), .R_WR(wRegEnTop_7_5), .R_In(wRegOut_7_5), .R_Out(wRegInTop_7_5) );
BHeap_Node #( 32 ) BHN_6_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_3), .P_In(wRegOut_6_3), .P_Out(wRegInBot_6_3), .L_WR(wRegEnTop_7_6), .L_In(wRegOut_7_6), .L_Out(wRegInTop_7_6), .R_WR(wRegEnTop_7_7), .R_In(wRegOut_7_7), .R_Out(wRegInTop_7_7) );
BHeap_Node #( 32 ) BHN_6_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_4), .P_In(wRegOut_6_4), .P_Out(wRegInBot_6_4), .L_WR(wRegEnTop_7_8), .L_In(wRegOut_7_8), .L_Out(wRegInTop_7_8), .R_WR(wRegEnTop_7_9), .R_In(wRegOut_7_9), .R_Out(wRegInTop_7_9) );
BHeap_Node #( 32 ) BHN_6_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_5), .P_In(wRegOut_6_5), .P_Out(wRegInBot_6_5), .L_WR(wRegEnTop_7_10), .L_In(wRegOut_7_10), .L_Out(wRegInTop_7_10), .R_WR(wRegEnTop_7_11), .R_In(wRegOut_7_11), .R_Out(wRegInTop_7_11) );
BHeap_Node #( 32 ) BHN_6_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_6), .P_In(wRegOut_6_6), .P_Out(wRegInBot_6_6), .L_WR(wRegEnTop_7_12), .L_In(wRegOut_7_12), .L_Out(wRegInTop_7_12), .R_WR(wRegEnTop_7_13), .R_In(wRegOut_7_13), .R_Out(wRegInTop_7_13) );
BHeap_Node #( 32 ) BHN_6_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_7), .P_In(wRegOut_6_7), .P_Out(wRegInBot_6_7), .L_WR(wRegEnTop_7_14), .L_In(wRegOut_7_14), .L_Out(wRegInTop_7_14), .R_WR(wRegEnTop_7_15), .R_In(wRegOut_7_15), .R_Out(wRegInTop_7_15) );
BHeap_Node #( 32 ) BHN_6_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_8), .P_In(wRegOut_6_8), .P_Out(wRegInBot_6_8), .L_WR(wRegEnTop_7_16), .L_In(wRegOut_7_16), .L_Out(wRegInTop_7_16), .R_WR(wRegEnTop_7_17), .R_In(wRegOut_7_17), .R_Out(wRegInTop_7_17) );
BHeap_Node #( 32 ) BHN_6_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_9), .P_In(wRegOut_6_9), .P_Out(wRegInBot_6_9), .L_WR(wRegEnTop_7_18), .L_In(wRegOut_7_18), .L_Out(wRegInTop_7_18), .R_WR(wRegEnTop_7_19), .R_In(wRegOut_7_19), .R_Out(wRegInTop_7_19) );
BHeap_Node #( 32 ) BHN_6_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_10), .P_In(wRegOut_6_10), .P_Out(wRegInBot_6_10), .L_WR(wRegEnTop_7_20), .L_In(wRegOut_7_20), .L_Out(wRegInTop_7_20), .R_WR(wRegEnTop_7_21), .R_In(wRegOut_7_21), .R_Out(wRegInTop_7_21) );
BHeap_Node #( 32 ) BHN_6_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_11), .P_In(wRegOut_6_11), .P_Out(wRegInBot_6_11), .L_WR(wRegEnTop_7_22), .L_In(wRegOut_7_22), .L_Out(wRegInTop_7_22), .R_WR(wRegEnTop_7_23), .R_In(wRegOut_7_23), .R_Out(wRegInTop_7_23) );
BHeap_Node #( 32 ) BHN_6_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_12), .P_In(wRegOut_6_12), .P_Out(wRegInBot_6_12), .L_WR(wRegEnTop_7_24), .L_In(wRegOut_7_24), .L_Out(wRegInTop_7_24), .R_WR(wRegEnTop_7_25), .R_In(wRegOut_7_25), .R_Out(wRegInTop_7_25) );
BHeap_Node #( 32 ) BHN_6_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_13), .P_In(wRegOut_6_13), .P_Out(wRegInBot_6_13), .L_WR(wRegEnTop_7_26), .L_In(wRegOut_7_26), .L_Out(wRegInTop_7_26), .R_WR(wRegEnTop_7_27), .R_In(wRegOut_7_27), .R_Out(wRegInTop_7_27) );
BHeap_Node #( 32 ) BHN_6_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_14), .P_In(wRegOut_6_14), .P_Out(wRegInBot_6_14), .L_WR(wRegEnTop_7_28), .L_In(wRegOut_7_28), .L_Out(wRegInTop_7_28), .R_WR(wRegEnTop_7_29), .R_In(wRegOut_7_29), .R_Out(wRegInTop_7_29) );
BHeap_Node #( 32 ) BHN_6_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_15), .P_In(wRegOut_6_15), .P_Out(wRegInBot_6_15), .L_WR(wRegEnTop_7_30), .L_In(wRegOut_7_30), .L_Out(wRegInTop_7_30), .R_WR(wRegEnTop_7_31), .R_In(wRegOut_7_31), .R_Out(wRegInTop_7_31) );
BHeap_Node #( 32 ) BHN_6_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_16), .P_In(wRegOut_6_16), .P_Out(wRegInBot_6_16), .L_WR(wRegEnTop_7_32), .L_In(wRegOut_7_32), .L_Out(wRegInTop_7_32), .R_WR(wRegEnTop_7_33), .R_In(wRegOut_7_33), .R_Out(wRegInTop_7_33) );
BHeap_Node #( 32 ) BHN_6_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_17), .P_In(wRegOut_6_17), .P_Out(wRegInBot_6_17), .L_WR(wRegEnTop_7_34), .L_In(wRegOut_7_34), .L_Out(wRegInTop_7_34), .R_WR(wRegEnTop_7_35), .R_In(wRegOut_7_35), .R_Out(wRegInTop_7_35) );
BHeap_Node #( 32 ) BHN_6_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_18), .P_In(wRegOut_6_18), .P_Out(wRegInBot_6_18), .L_WR(wRegEnTop_7_36), .L_In(wRegOut_7_36), .L_Out(wRegInTop_7_36), .R_WR(wRegEnTop_7_37), .R_In(wRegOut_7_37), .R_Out(wRegInTop_7_37) );
BHeap_Node #( 32 ) BHN_6_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_19), .P_In(wRegOut_6_19), .P_Out(wRegInBot_6_19), .L_WR(wRegEnTop_7_38), .L_In(wRegOut_7_38), .L_Out(wRegInTop_7_38), .R_WR(wRegEnTop_7_39), .R_In(wRegOut_7_39), .R_Out(wRegInTop_7_39) );
BHeap_Node #( 32 ) BHN_6_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_20), .P_In(wRegOut_6_20), .P_Out(wRegInBot_6_20), .L_WR(wRegEnTop_7_40), .L_In(wRegOut_7_40), .L_Out(wRegInTop_7_40), .R_WR(wRegEnTop_7_41), .R_In(wRegOut_7_41), .R_Out(wRegInTop_7_41) );
BHeap_Node #( 32 ) BHN_6_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_21), .P_In(wRegOut_6_21), .P_Out(wRegInBot_6_21), .L_WR(wRegEnTop_7_42), .L_In(wRegOut_7_42), .L_Out(wRegInTop_7_42), .R_WR(wRegEnTop_7_43), .R_In(wRegOut_7_43), .R_Out(wRegInTop_7_43) );
BHeap_Node #( 32 ) BHN_6_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_22), .P_In(wRegOut_6_22), .P_Out(wRegInBot_6_22), .L_WR(wRegEnTop_7_44), .L_In(wRegOut_7_44), .L_Out(wRegInTop_7_44), .R_WR(wRegEnTop_7_45), .R_In(wRegOut_7_45), .R_Out(wRegInTop_7_45) );
BHeap_Node #( 32 ) BHN_6_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_23), .P_In(wRegOut_6_23), .P_Out(wRegInBot_6_23), .L_WR(wRegEnTop_7_46), .L_In(wRegOut_7_46), .L_Out(wRegInTop_7_46), .R_WR(wRegEnTop_7_47), .R_In(wRegOut_7_47), .R_Out(wRegInTop_7_47) );
BHeap_Node #( 32 ) BHN_6_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_24), .P_In(wRegOut_6_24), .P_Out(wRegInBot_6_24), .L_WR(wRegEnTop_7_48), .L_In(wRegOut_7_48), .L_Out(wRegInTop_7_48), .R_WR(wRegEnTop_7_49), .R_In(wRegOut_7_49), .R_Out(wRegInTop_7_49) );
BHeap_Node #( 32 ) BHN_6_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_25), .P_In(wRegOut_6_25), .P_Out(wRegInBot_6_25), .L_WR(wRegEnTop_7_50), .L_In(wRegOut_7_50), .L_Out(wRegInTop_7_50), .R_WR(wRegEnTop_7_51), .R_In(wRegOut_7_51), .R_Out(wRegInTop_7_51) );
BHeap_Node #( 32 ) BHN_6_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_26), .P_In(wRegOut_6_26), .P_Out(wRegInBot_6_26), .L_WR(wRegEnTop_7_52), .L_In(wRegOut_7_52), .L_Out(wRegInTop_7_52), .R_WR(wRegEnTop_7_53), .R_In(wRegOut_7_53), .R_Out(wRegInTop_7_53) );
BHeap_Node #( 32 ) BHN_6_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_27), .P_In(wRegOut_6_27), .P_Out(wRegInBot_6_27), .L_WR(wRegEnTop_7_54), .L_In(wRegOut_7_54), .L_Out(wRegInTop_7_54), .R_WR(wRegEnTop_7_55), .R_In(wRegOut_7_55), .R_Out(wRegInTop_7_55) );
BHeap_Node #( 32 ) BHN_6_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_28), .P_In(wRegOut_6_28), .P_Out(wRegInBot_6_28), .L_WR(wRegEnTop_7_56), .L_In(wRegOut_7_56), .L_Out(wRegInTop_7_56), .R_WR(wRegEnTop_7_57), .R_In(wRegOut_7_57), .R_Out(wRegInTop_7_57) );
BHeap_Node #( 32 ) BHN_6_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_29), .P_In(wRegOut_6_29), .P_Out(wRegInBot_6_29), .L_WR(wRegEnTop_7_58), .L_In(wRegOut_7_58), .L_Out(wRegInTop_7_58), .R_WR(wRegEnTop_7_59), .R_In(wRegOut_7_59), .R_Out(wRegInTop_7_59) );
BHeap_Node #( 32 ) BHN_6_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_30), .P_In(wRegOut_6_30), .P_Out(wRegInBot_6_30), .L_WR(wRegEnTop_7_60), .L_In(wRegOut_7_60), .L_Out(wRegInTop_7_60), .R_WR(wRegEnTop_7_61), .R_In(wRegOut_7_61), .R_Out(wRegInTop_7_61) );
BHeap_Node #( 32 ) BHN_6_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_31), .P_In(wRegOut_6_31), .P_Out(wRegInBot_6_31), .L_WR(wRegEnTop_7_62), .L_In(wRegOut_7_62), .L_Out(wRegInTop_7_62), .R_WR(wRegEnTop_7_63), .R_In(wRegOut_7_63), .R_Out(wRegInTop_7_63) );
BHeap_Node #( 32 ) BHN_6_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_32), .P_In(wRegOut_6_32), .P_Out(wRegInBot_6_32), .L_WR(wRegEnTop_7_64), .L_In(wRegOut_7_64), .L_Out(wRegInTop_7_64), .R_WR(wRegEnTop_7_65), .R_In(wRegOut_7_65), .R_Out(wRegInTop_7_65) );
BHeap_Node #( 32 ) BHN_6_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_33), .P_In(wRegOut_6_33), .P_Out(wRegInBot_6_33), .L_WR(wRegEnTop_7_66), .L_In(wRegOut_7_66), .L_Out(wRegInTop_7_66), .R_WR(wRegEnTop_7_67), .R_In(wRegOut_7_67), .R_Out(wRegInTop_7_67) );
BHeap_Node #( 32 ) BHN_6_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_34), .P_In(wRegOut_6_34), .P_Out(wRegInBot_6_34), .L_WR(wRegEnTop_7_68), .L_In(wRegOut_7_68), .L_Out(wRegInTop_7_68), .R_WR(wRegEnTop_7_69), .R_In(wRegOut_7_69), .R_Out(wRegInTop_7_69) );
BHeap_Node #( 32 ) BHN_6_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_35), .P_In(wRegOut_6_35), .P_Out(wRegInBot_6_35), .L_WR(wRegEnTop_7_70), .L_In(wRegOut_7_70), .L_Out(wRegInTop_7_70), .R_WR(wRegEnTop_7_71), .R_In(wRegOut_7_71), .R_Out(wRegInTop_7_71) );
BHeap_Node #( 32 ) BHN_6_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_36), .P_In(wRegOut_6_36), .P_Out(wRegInBot_6_36), .L_WR(wRegEnTop_7_72), .L_In(wRegOut_7_72), .L_Out(wRegInTop_7_72), .R_WR(wRegEnTop_7_73), .R_In(wRegOut_7_73), .R_Out(wRegInTop_7_73) );
BHeap_Node #( 32 ) BHN_6_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_37), .P_In(wRegOut_6_37), .P_Out(wRegInBot_6_37), .L_WR(wRegEnTop_7_74), .L_In(wRegOut_7_74), .L_Out(wRegInTop_7_74), .R_WR(wRegEnTop_7_75), .R_In(wRegOut_7_75), .R_Out(wRegInTop_7_75) );
BHeap_Node #( 32 ) BHN_6_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_38), .P_In(wRegOut_6_38), .P_Out(wRegInBot_6_38), .L_WR(wRegEnTop_7_76), .L_In(wRegOut_7_76), .L_Out(wRegInTop_7_76), .R_WR(wRegEnTop_7_77), .R_In(wRegOut_7_77), .R_Out(wRegInTop_7_77) );
BHeap_Node #( 32 ) BHN_6_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_39), .P_In(wRegOut_6_39), .P_Out(wRegInBot_6_39), .L_WR(wRegEnTop_7_78), .L_In(wRegOut_7_78), .L_Out(wRegInTop_7_78), .R_WR(wRegEnTop_7_79), .R_In(wRegOut_7_79), .R_Out(wRegInTop_7_79) );
BHeap_Node #( 32 ) BHN_6_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_40), .P_In(wRegOut_6_40), .P_Out(wRegInBot_6_40), .L_WR(wRegEnTop_7_80), .L_In(wRegOut_7_80), .L_Out(wRegInTop_7_80), .R_WR(wRegEnTop_7_81), .R_In(wRegOut_7_81), .R_Out(wRegInTop_7_81) );
BHeap_Node #( 32 ) BHN_6_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_41), .P_In(wRegOut_6_41), .P_Out(wRegInBot_6_41), .L_WR(wRegEnTop_7_82), .L_In(wRegOut_7_82), .L_Out(wRegInTop_7_82), .R_WR(wRegEnTop_7_83), .R_In(wRegOut_7_83), .R_Out(wRegInTop_7_83) );
BHeap_Node #( 32 ) BHN_6_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_42), .P_In(wRegOut_6_42), .P_Out(wRegInBot_6_42), .L_WR(wRegEnTop_7_84), .L_In(wRegOut_7_84), .L_Out(wRegInTop_7_84), .R_WR(wRegEnTop_7_85), .R_In(wRegOut_7_85), .R_Out(wRegInTop_7_85) );
BHeap_Node #( 32 ) BHN_6_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_43), .P_In(wRegOut_6_43), .P_Out(wRegInBot_6_43), .L_WR(wRegEnTop_7_86), .L_In(wRegOut_7_86), .L_Out(wRegInTop_7_86), .R_WR(wRegEnTop_7_87), .R_In(wRegOut_7_87), .R_Out(wRegInTop_7_87) );
BHeap_Node #( 32 ) BHN_6_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_44), .P_In(wRegOut_6_44), .P_Out(wRegInBot_6_44), .L_WR(wRegEnTop_7_88), .L_In(wRegOut_7_88), .L_Out(wRegInTop_7_88), .R_WR(wRegEnTop_7_89), .R_In(wRegOut_7_89), .R_Out(wRegInTop_7_89) );
BHeap_Node #( 32 ) BHN_6_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_45), .P_In(wRegOut_6_45), .P_Out(wRegInBot_6_45), .L_WR(wRegEnTop_7_90), .L_In(wRegOut_7_90), .L_Out(wRegInTop_7_90), .R_WR(wRegEnTop_7_91), .R_In(wRegOut_7_91), .R_Out(wRegInTop_7_91) );
BHeap_Node #( 32 ) BHN_6_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_46), .P_In(wRegOut_6_46), .P_Out(wRegInBot_6_46), .L_WR(wRegEnTop_7_92), .L_In(wRegOut_7_92), .L_Out(wRegInTop_7_92), .R_WR(wRegEnTop_7_93), .R_In(wRegOut_7_93), .R_Out(wRegInTop_7_93) );
BHeap_Node #( 32 ) BHN_6_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_47), .P_In(wRegOut_6_47), .P_Out(wRegInBot_6_47), .L_WR(wRegEnTop_7_94), .L_In(wRegOut_7_94), .L_Out(wRegInTop_7_94), .R_WR(wRegEnTop_7_95), .R_In(wRegOut_7_95), .R_Out(wRegInTop_7_95) );
BHeap_Node #( 32 ) BHN_6_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_48), .P_In(wRegOut_6_48), .P_Out(wRegInBot_6_48), .L_WR(wRegEnTop_7_96), .L_In(wRegOut_7_96), .L_Out(wRegInTop_7_96), .R_WR(wRegEnTop_7_97), .R_In(wRegOut_7_97), .R_Out(wRegInTop_7_97) );
BHeap_Node #( 32 ) BHN_6_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_49), .P_In(wRegOut_6_49), .P_Out(wRegInBot_6_49), .L_WR(wRegEnTop_7_98), .L_In(wRegOut_7_98), .L_Out(wRegInTop_7_98), .R_WR(wRegEnTop_7_99), .R_In(wRegOut_7_99), .R_Out(wRegInTop_7_99) );
BHeap_Node #( 32 ) BHN_6_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_50), .P_In(wRegOut_6_50), .P_Out(wRegInBot_6_50), .L_WR(wRegEnTop_7_100), .L_In(wRegOut_7_100), .L_Out(wRegInTop_7_100), .R_WR(wRegEnTop_7_101), .R_In(wRegOut_7_101), .R_Out(wRegInTop_7_101) );
BHeap_Node #( 32 ) BHN_6_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_51), .P_In(wRegOut_6_51), .P_Out(wRegInBot_6_51), .L_WR(wRegEnTop_7_102), .L_In(wRegOut_7_102), .L_Out(wRegInTop_7_102), .R_WR(wRegEnTop_7_103), .R_In(wRegOut_7_103), .R_Out(wRegInTop_7_103) );
BHeap_Node #( 32 ) BHN_6_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_52), .P_In(wRegOut_6_52), .P_Out(wRegInBot_6_52), .L_WR(wRegEnTop_7_104), .L_In(wRegOut_7_104), .L_Out(wRegInTop_7_104), .R_WR(wRegEnTop_7_105), .R_In(wRegOut_7_105), .R_Out(wRegInTop_7_105) );
BHeap_Node #( 32 ) BHN_6_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_53), .P_In(wRegOut_6_53), .P_Out(wRegInBot_6_53), .L_WR(wRegEnTop_7_106), .L_In(wRegOut_7_106), .L_Out(wRegInTop_7_106), .R_WR(wRegEnTop_7_107), .R_In(wRegOut_7_107), .R_Out(wRegInTop_7_107) );
BHeap_Node #( 32 ) BHN_6_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_54), .P_In(wRegOut_6_54), .P_Out(wRegInBot_6_54), .L_WR(wRegEnTop_7_108), .L_In(wRegOut_7_108), .L_Out(wRegInTop_7_108), .R_WR(wRegEnTop_7_109), .R_In(wRegOut_7_109), .R_Out(wRegInTop_7_109) );
BHeap_Node #( 32 ) BHN_6_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_55), .P_In(wRegOut_6_55), .P_Out(wRegInBot_6_55), .L_WR(wRegEnTop_7_110), .L_In(wRegOut_7_110), .L_Out(wRegInTop_7_110), .R_WR(wRegEnTop_7_111), .R_In(wRegOut_7_111), .R_Out(wRegInTop_7_111) );
BHeap_Node #( 32 ) BHN_6_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_56), .P_In(wRegOut_6_56), .P_Out(wRegInBot_6_56), .L_WR(wRegEnTop_7_112), .L_In(wRegOut_7_112), .L_Out(wRegInTop_7_112), .R_WR(wRegEnTop_7_113), .R_In(wRegOut_7_113), .R_Out(wRegInTop_7_113) );
BHeap_Node #( 32 ) BHN_6_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_57), .P_In(wRegOut_6_57), .P_Out(wRegInBot_6_57), .L_WR(wRegEnTop_7_114), .L_In(wRegOut_7_114), .L_Out(wRegInTop_7_114), .R_WR(wRegEnTop_7_115), .R_In(wRegOut_7_115), .R_Out(wRegInTop_7_115) );
BHeap_Node #( 32 ) BHN_6_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_58), .P_In(wRegOut_6_58), .P_Out(wRegInBot_6_58), .L_WR(wRegEnTop_7_116), .L_In(wRegOut_7_116), .L_Out(wRegInTop_7_116), .R_WR(wRegEnTop_7_117), .R_In(wRegOut_7_117), .R_Out(wRegInTop_7_117) );
BHeap_Node #( 32 ) BHN_6_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_59), .P_In(wRegOut_6_59), .P_Out(wRegInBot_6_59), .L_WR(wRegEnTop_7_118), .L_In(wRegOut_7_118), .L_Out(wRegInTop_7_118), .R_WR(wRegEnTop_7_119), .R_In(wRegOut_7_119), .R_Out(wRegInTop_7_119) );
BHeap_Node #( 32 ) BHN_6_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_60), .P_In(wRegOut_6_60), .P_Out(wRegInBot_6_60), .L_WR(wRegEnTop_7_120), .L_In(wRegOut_7_120), .L_Out(wRegInTop_7_120), .R_WR(wRegEnTop_7_121), .R_In(wRegOut_7_121), .R_Out(wRegInTop_7_121) );
BHeap_Node #( 32 ) BHN_6_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_61), .P_In(wRegOut_6_61), .P_Out(wRegInBot_6_61), .L_WR(wRegEnTop_7_122), .L_In(wRegOut_7_122), .L_Out(wRegInTop_7_122), .R_WR(wRegEnTop_7_123), .R_In(wRegOut_7_123), .R_Out(wRegInTop_7_123) );
BHeap_Node #( 32 ) BHN_6_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_62), .P_In(wRegOut_6_62), .P_Out(wRegInBot_6_62), .L_WR(wRegEnTop_7_124), .L_In(wRegOut_7_124), .L_Out(wRegInTop_7_124), .R_WR(wRegEnTop_7_125), .R_In(wRegOut_7_125), .R_Out(wRegInTop_7_125) );
BHeap_Node #( 32 ) BHN_6_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Enable(wEnable_6), .P_WR(wRegEnBot_6_63), .P_In(wRegOut_6_63), .P_Out(wRegInBot_6_63), .L_WR(wRegEnTop_7_126), .L_In(wRegOut_7_126), .L_Out(wRegInTop_7_126), .R_WR(wRegEnTop_7_127), .R_In(wRegOut_7_127), .R_Out(wRegInTop_7_127) );
BHeap_CtrlReg #( 32 ) BHCR_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_1), .Out(wCtrlOut_0), .Enable(wEnable_0) );
BHeap_CtrlReg #( 32 ) BHCR_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_2), .Out(wCtrlOut_1), .Enable(wEnable_1) );
BHeap_CtrlReg #( 32 ) BHCR_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_3), .Out(wCtrlOut_2), .Enable(wEnable_2) );
BHeap_CtrlReg #( 32 ) BHCR_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_4), .Out(wCtrlOut_3), .Enable(wEnable_3) );
BHeap_CtrlReg #( 32 ) BHCR_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_5), .Out(wCtrlOut_4), .Enable(wEnable_4) );
BHeap_CtrlReg #( 32 ) BHCR_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_6), .Out(wCtrlOut_5), .Enable(wEnable_5) );
BHeap_CtrlReg #( 32 ) BHCR_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .In(wCtrlOut_7), .Out(wCtrlOut_6), .Enable(wEnable_6) );
BHeap_Control #( 4, 1, 32, 1 ) BHC ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Go(wCtrlOut_7), .Done(wCtrlOut_0), .ScanIn(ScanLink0), .ScanOut(ScanLink255), .ScanEnable(ScanEnable), .ScanId(1'd0) );

/*
 *
 * RAW Benchmark Suite main module trailer
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
