

/*
 *
 * RAW Benchmark Suite main defines
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz 

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/jacobi/src/library.v,v 1.5 1997/08/09 05:57:41 jbabb Exp $
 *
 * Library for Jacobi benchmark
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 * This is the behavioral verilog library for this benchmark.
 * By convention, all module names start with the benchmark name.
 * All top-level modules must have the global connections:
 *   Clk, Reset, RD, WR, Addr, DataIn, DataOut
 * Modules may also have any number of local connections or
 * sub-modules without restriction.
 *
 */


/* The basic array node */

module Jacobi_Node (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		    ScanIn, ScanOut, ScanEnable,
		    Id, Enable, NorthIn, SouthIn, EastIn, WestIn, Out);
   
   parameter WIDTH    = 8,
	     IDWIDTH  = 8,
	     BOUNDARY = 0,
	     SCAN     = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;   


   /* local connections */
   
   input			 Enable;
   input [IDWIDTH-1:0]		 Id;
   input [WIDTH-1:0]		 NorthIn,SouthIn,EastIn,WestIn;
   output [WIDTH-1:0]		 Out;
   
   reg [WIDTH-1:0]		 Out;
   
   
   /* support reading of the node data value (non-scan only) */
   
   assign DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out: `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;

   
   always @(posedge Clk)
      begin	

	 
	 /* reset will initialize the entire array to zero */
	 
	 if (Reset)
	    Out=0;	 


	 /* support scan in */

	 else if (SCAN && ScanEnable)
	    Out=ScanIn[WIDTH-1:0];
	 

	 /* support writing of the node data value (non-scan only) */
	 
	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0]==Id))
	    Out=DataIn[WIDTH-1:0];
	 

	 /* for non-boundary nodes, do the Jacobi computation when enabled */
	 
	 else if (!BOUNDARY && Enable)
	    Out=(NorthIn+SouthIn+EastIn+WestIn) >> 2;

      end
endmodule


/* 
 * A control module to count iterations.
 *
 * Writing to Address==ID will set a counter.
 *
 * The other Jacobi nodes will be enabled by this module when 
 * count is greater than zero.
 *
 * The counter will decrement every cycle down to zero.
 *
 * This module also handles scan control.
 */

module Jacobi_Control (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		       ScanIn, ScanOut, ScanEnable,
		       Id,ScanId,Enable);
   
   parameter WIDTH   = 8,
	     CWIDTH  = 8,
	     IDWIDTH = 8,
	     SCAN    = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [IDWIDTH-1:0]		 ScanId;
   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;   


   /* local connections */
   
   input [IDWIDTH-1:0]		 Id;
   output			 Enable;
   
   
   /* a register for the counter and scan */

   reg [CWIDTH-1:0]		 count;
   reg [WIDTH-1:0]		 ScanReg;

   
   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? count:
      (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;
   
   
   /* enable when count is active */
   
   assign Enable = !(count==0);

   
   always @(posedge Clk)
      begin

	 
	 /* store current scan output */

	 ScanReg=ScanIn;


	 /* Logic to reset, write, and decrement the counter */
	 
	 if (Reset)
	    count=0;
	 else if (WR && (Addr[IDWIDTH-1:0]==Id))
	    count=DataIn[CWIDTH-1:0];
	 else if(count) 
	    count=count-1;
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [7:0] nOut0_0;
wire [7:0] nScanOut0;
wire [7:0] nOut0_1;
wire [7:0] nScanOut1;
wire [7:0] nOut0_2;
wire [7:0] nScanOut2;
wire [7:0] nOut0_3;
wire [7:0] nScanOut3;
wire [7:0] nOut0_4;
wire [7:0] nScanOut4;
wire [7:0] nOut0_5;
wire [7:0] nScanOut5;
wire [7:0] nOut0_6;
wire [7:0] nScanOut6;
wire [7:0] nOut0_7;
wire [7:0] nScanOut7;
wire [7:0] nOut0_8;
wire [7:0] nScanOut8;
wire [7:0] nOut0_9;
wire [7:0] nScanOut9;
wire [7:0] nOut0_10;
wire [7:0] nScanOut10;
wire [7:0] nOut0_11;
wire [7:0] nScanOut11;
wire [7:0] nOut0_12;
wire [7:0] nScanOut12;
wire [7:0] nOut0_13;
wire [7:0] nScanOut13;
wire [7:0] nOut0_14;
wire [7:0] nScanOut14;
wire [7:0] nOut0_15;
wire [7:0] nScanOut15;
wire [7:0] nOut1_0;
wire [7:0] nScanOut16;
wire [7:0] nOut1_1;
wire [7:0] nScanOut17;
wire [7:0] nOut1_2;
wire [7:0] nScanOut18;
wire [7:0] nOut1_3;
wire [7:0] nScanOut19;
wire [7:0] nOut1_4;
wire [7:0] nScanOut20;
wire [7:0] nOut1_5;
wire [7:0] nScanOut21;
wire [7:0] nOut1_6;
wire [7:0] nScanOut22;
wire [7:0] nOut1_7;
wire [7:0] nScanOut23;
wire [7:0] nOut1_8;
wire [7:0] nScanOut24;
wire [7:0] nOut1_9;
wire [7:0] nScanOut25;
wire [7:0] nOut1_10;
wire [7:0] nScanOut26;
wire [7:0] nOut1_11;
wire [7:0] nScanOut27;
wire [7:0] nOut1_12;
wire [7:0] nScanOut28;
wire [7:0] nOut1_13;
wire [7:0] nScanOut29;
wire [7:0] nOut1_14;
wire [7:0] nScanOut30;
wire [7:0] nOut1_15;
wire [7:0] nScanOut31;
wire [7:0] nOut2_0;
wire [7:0] nScanOut32;
wire [7:0] nOut2_1;
wire [7:0] nScanOut33;
wire [7:0] nOut2_2;
wire [7:0] nScanOut34;
wire [7:0] nOut2_3;
wire [7:0] nScanOut35;
wire [7:0] nOut2_4;
wire [7:0] nScanOut36;
wire [7:0] nOut2_5;
wire [7:0] nScanOut37;
wire [7:0] nOut2_6;
wire [7:0] nScanOut38;
wire [7:0] nOut2_7;
wire [7:0] nScanOut39;
wire [7:0] nOut2_8;
wire [7:0] nScanOut40;
wire [7:0] nOut2_9;
wire [7:0] nScanOut41;
wire [7:0] nOut2_10;
wire [7:0] nScanOut42;
wire [7:0] nOut2_11;
wire [7:0] nScanOut43;
wire [7:0] nOut2_12;
wire [7:0] nScanOut44;
wire [7:0] nOut2_13;
wire [7:0] nScanOut45;
wire [7:0] nOut2_14;
wire [7:0] nScanOut46;
wire [7:0] nOut2_15;
wire [7:0] nScanOut47;
wire [7:0] nOut3_0;
wire [7:0] nScanOut48;
wire [7:0] nOut3_1;
wire [7:0] nScanOut49;
wire [7:0] nOut3_2;
wire [7:0] nScanOut50;
wire [7:0] nOut3_3;
wire [7:0] nScanOut51;
wire [7:0] nOut3_4;
wire [7:0] nScanOut52;
wire [7:0] nOut3_5;
wire [7:0] nScanOut53;
wire [7:0] nOut3_6;
wire [7:0] nScanOut54;
wire [7:0] nOut3_7;
wire [7:0] nScanOut55;
wire [7:0] nOut3_8;
wire [7:0] nScanOut56;
wire [7:0] nOut3_9;
wire [7:0] nScanOut57;
wire [7:0] nOut3_10;
wire [7:0] nScanOut58;
wire [7:0] nOut3_11;
wire [7:0] nScanOut59;
wire [7:0] nOut3_12;
wire [7:0] nScanOut60;
wire [7:0] nOut3_13;
wire [7:0] nScanOut61;
wire [7:0] nOut3_14;
wire [7:0] nScanOut62;
wire [7:0] nOut3_15;
wire [7:0] nScanOut63;
wire [7:0] nOut4_0;
wire [7:0] nScanOut64;
wire [7:0] nOut4_1;
wire [7:0] nScanOut65;
wire [7:0] nOut4_2;
wire [7:0] nScanOut66;
wire [7:0] nOut4_3;
wire [7:0] nScanOut67;
wire [7:0] nOut4_4;
wire [7:0] nScanOut68;
wire [7:0] nOut4_5;
wire [7:0] nScanOut69;
wire [7:0] nOut4_6;
wire [7:0] nScanOut70;
wire [7:0] nOut4_7;
wire [7:0] nScanOut71;
wire [7:0] nOut4_8;
wire [7:0] nScanOut72;
wire [7:0] nOut4_9;
wire [7:0] nScanOut73;
wire [7:0] nOut4_10;
wire [7:0] nScanOut74;
wire [7:0] nOut4_11;
wire [7:0] nScanOut75;
wire [7:0] nOut4_12;
wire [7:0] nScanOut76;
wire [7:0] nOut4_13;
wire [7:0] nScanOut77;
wire [7:0] nOut4_14;
wire [7:0] nScanOut78;
wire [7:0] nOut4_15;
wire [7:0] nScanOut79;
wire [7:0] nOut5_0;
wire [7:0] nScanOut80;
wire [7:0] nOut5_1;
wire [7:0] nScanOut81;
wire [7:0] nOut5_2;
wire [7:0] nScanOut82;
wire [7:0] nOut5_3;
wire [7:0] nScanOut83;
wire [7:0] nOut5_4;
wire [7:0] nScanOut84;
wire [7:0] nOut5_5;
wire [7:0] nScanOut85;
wire [7:0] nOut5_6;
wire [7:0] nScanOut86;
wire [7:0] nOut5_7;
wire [7:0] nScanOut87;
wire [7:0] nOut5_8;
wire [7:0] nScanOut88;
wire [7:0] nOut5_9;
wire [7:0] nScanOut89;
wire [7:0] nOut5_10;
wire [7:0] nScanOut90;
wire [7:0] nOut5_11;
wire [7:0] nScanOut91;
wire [7:0] nOut5_12;
wire [7:0] nScanOut92;
wire [7:0] nOut5_13;
wire [7:0] nScanOut93;
wire [7:0] nOut5_14;
wire [7:0] nScanOut94;
wire [7:0] nOut5_15;
wire [7:0] nScanOut95;
wire [7:0] nOut6_0;
wire [7:0] nScanOut96;
wire [7:0] nOut6_1;
wire [7:0] nScanOut97;
wire [7:0] nOut6_2;
wire [7:0] nScanOut98;
wire [7:0] nOut6_3;
wire [7:0] nScanOut99;
wire [7:0] nOut6_4;
wire [7:0] nScanOut100;
wire [7:0] nOut6_5;
wire [7:0] nScanOut101;
wire [7:0] nOut6_6;
wire [7:0] nScanOut102;
wire [7:0] nOut6_7;
wire [7:0] nScanOut103;
wire [7:0] nOut6_8;
wire [7:0] nScanOut104;
wire [7:0] nOut6_9;
wire [7:0] nScanOut105;
wire [7:0] nOut6_10;
wire [7:0] nScanOut106;
wire [7:0] nOut6_11;
wire [7:0] nScanOut107;
wire [7:0] nOut6_12;
wire [7:0] nScanOut108;
wire [7:0] nOut6_13;
wire [7:0] nScanOut109;
wire [7:0] nOut6_14;
wire [7:0] nScanOut110;
wire [7:0] nOut6_15;
wire [7:0] nScanOut111;
wire [7:0] nOut7_0;
wire [7:0] nScanOut112;
wire [7:0] nOut7_1;
wire [7:0] nScanOut113;
wire [7:0] nOut7_2;
wire [7:0] nScanOut114;
wire [7:0] nOut7_3;
wire [7:0] nScanOut115;
wire [7:0] nOut7_4;
wire [7:0] nScanOut116;
wire [7:0] nOut7_5;
wire [7:0] nScanOut117;
wire [7:0] nOut7_6;
wire [7:0] nScanOut118;
wire [7:0] nOut7_7;
wire [7:0] nScanOut119;
wire [7:0] nOut7_8;
wire [7:0] nScanOut120;
wire [7:0] nOut7_9;
wire [7:0] nScanOut121;
wire [7:0] nOut7_10;
wire [7:0] nScanOut122;
wire [7:0] nOut7_11;
wire [7:0] nScanOut123;
wire [7:0] nOut7_12;
wire [7:0] nScanOut124;
wire [7:0] nOut7_13;
wire [7:0] nScanOut125;
wire [7:0] nOut7_14;
wire [7:0] nScanOut126;
wire [7:0] nOut7_15;
wire [7:0] nScanOut127;
wire [7:0] nOut8_0;
wire [7:0] nScanOut128;
wire [7:0] nOut8_1;
wire [7:0] nScanOut129;
wire [7:0] nOut8_2;
wire [7:0] nScanOut130;
wire [7:0] nOut8_3;
wire [7:0] nScanOut131;
wire [7:0] nOut8_4;
wire [7:0] nScanOut132;
wire [7:0] nOut8_5;
wire [7:0] nScanOut133;
wire [7:0] nOut8_6;
wire [7:0] nScanOut134;
wire [7:0] nOut8_7;
wire [7:0] nScanOut135;
wire [7:0] nOut8_8;
wire [7:0] nScanOut136;
wire [7:0] nOut8_9;
wire [7:0] nScanOut137;
wire [7:0] nOut8_10;
wire [7:0] nScanOut138;
wire [7:0] nOut8_11;
wire [7:0] nScanOut139;
wire [7:0] nOut8_12;
wire [7:0] nScanOut140;
wire [7:0] nOut8_13;
wire [7:0] nScanOut141;
wire [7:0] nOut8_14;
wire [7:0] nScanOut142;
wire [7:0] nOut8_15;
wire [7:0] nScanOut143;
wire [7:0] nOut9_0;
wire [7:0] nScanOut144;
wire [7:0] nOut9_1;
wire [7:0] nScanOut145;
wire [7:0] nOut9_2;
wire [7:0] nScanOut146;
wire [7:0] nOut9_3;
wire [7:0] nScanOut147;
wire [7:0] nOut9_4;
wire [7:0] nScanOut148;
wire [7:0] nOut9_5;
wire [7:0] nScanOut149;
wire [7:0] nOut9_6;
wire [7:0] nScanOut150;
wire [7:0] nOut9_7;
wire [7:0] nScanOut151;
wire [7:0] nOut9_8;
wire [7:0] nScanOut152;
wire [7:0] nOut9_9;
wire [7:0] nScanOut153;
wire [7:0] nOut9_10;
wire [7:0] nScanOut154;
wire [7:0] nOut9_11;
wire [7:0] nScanOut155;
wire [7:0] nOut9_12;
wire [7:0] nScanOut156;
wire [7:0] nOut9_13;
wire [7:0] nScanOut157;
wire [7:0] nOut9_14;
wire [7:0] nScanOut158;
wire [7:0] nOut9_15;
wire [7:0] nScanOut159;
wire [7:0] nOut10_0;
wire [7:0] nScanOut160;
wire [7:0] nOut10_1;
wire [7:0] nScanOut161;
wire [7:0] nOut10_2;
wire [7:0] nScanOut162;
wire [7:0] nOut10_3;
wire [7:0] nScanOut163;
wire [7:0] nOut10_4;
wire [7:0] nScanOut164;
wire [7:0] nOut10_5;
wire [7:0] nScanOut165;
wire [7:0] nOut10_6;
wire [7:0] nScanOut166;
wire [7:0] nOut10_7;
wire [7:0] nScanOut167;
wire [7:0] nOut10_8;
wire [7:0] nScanOut168;
wire [7:0] nOut10_9;
wire [7:0] nScanOut169;
wire [7:0] nOut10_10;
wire [7:0] nScanOut170;
wire [7:0] nOut10_11;
wire [7:0] nScanOut171;
wire [7:0] nOut10_12;
wire [7:0] nScanOut172;
wire [7:0] nOut10_13;
wire [7:0] nScanOut173;
wire [7:0] nOut10_14;
wire [7:0] nScanOut174;
wire [7:0] nOut10_15;
wire [7:0] nScanOut175;
wire [7:0] nOut11_0;
wire [7:0] nScanOut176;
wire [7:0] nOut11_1;
wire [7:0] nScanOut177;
wire [7:0] nOut11_2;
wire [7:0] nScanOut178;
wire [7:0] nOut11_3;
wire [7:0] nScanOut179;
wire [7:0] nOut11_4;
wire [7:0] nScanOut180;
wire [7:0] nOut11_5;
wire [7:0] nScanOut181;
wire [7:0] nOut11_6;
wire [7:0] nScanOut182;
wire [7:0] nOut11_7;
wire [7:0] nScanOut183;
wire [7:0] nOut11_8;
wire [7:0] nScanOut184;
wire [7:0] nOut11_9;
wire [7:0] nScanOut185;
wire [7:0] nOut11_10;
wire [7:0] nScanOut186;
wire [7:0] nOut11_11;
wire [7:0] nScanOut187;
wire [7:0] nOut11_12;
wire [7:0] nScanOut188;
wire [7:0] nOut11_13;
wire [7:0] nScanOut189;
wire [7:0] nOut11_14;
wire [7:0] nScanOut190;
wire [7:0] nOut11_15;
wire [7:0] nScanOut191;
wire [7:0] nOut12_0;
wire [7:0] nScanOut192;
wire [7:0] nOut12_1;
wire [7:0] nScanOut193;
wire [7:0] nOut12_2;
wire [7:0] nScanOut194;
wire [7:0] nOut12_3;
wire [7:0] nScanOut195;
wire [7:0] nOut12_4;
wire [7:0] nScanOut196;
wire [7:0] nOut12_5;
wire [7:0] nScanOut197;
wire [7:0] nOut12_6;
wire [7:0] nScanOut198;
wire [7:0] nOut12_7;
wire [7:0] nScanOut199;
wire [7:0] nOut12_8;
wire [7:0] nScanOut200;
wire [7:0] nOut12_9;
wire [7:0] nScanOut201;
wire [7:0] nOut12_10;
wire [7:0] nScanOut202;
wire [7:0] nOut12_11;
wire [7:0] nScanOut203;
wire [7:0] nOut12_12;
wire [7:0] nScanOut204;
wire [7:0] nOut12_13;
wire [7:0] nScanOut205;
wire [7:0] nOut12_14;
wire [7:0] nScanOut206;
wire [7:0] nOut12_15;
wire [7:0] nScanOut207;
wire [7:0] nOut13_0;
wire [7:0] nScanOut208;
wire [7:0] nOut13_1;
wire [7:0] nScanOut209;
wire [7:0] nOut13_2;
wire [7:0] nScanOut210;
wire [7:0] nOut13_3;
wire [7:0] nScanOut211;
wire [7:0] nOut13_4;
wire [7:0] nScanOut212;
wire [7:0] nOut13_5;
wire [7:0] nScanOut213;
wire [7:0] nOut13_6;
wire [7:0] nScanOut214;
wire [7:0] nOut13_7;
wire [7:0] nScanOut215;
wire [7:0] nOut13_8;
wire [7:0] nScanOut216;
wire [7:0] nOut13_9;
wire [7:0] nScanOut217;
wire [7:0] nOut13_10;
wire [7:0] nScanOut218;
wire [7:0] nOut13_11;
wire [7:0] nScanOut219;
wire [7:0] nOut13_12;
wire [7:0] nScanOut220;
wire [7:0] nOut13_13;
wire [7:0] nScanOut221;
wire [7:0] nOut13_14;
wire [7:0] nScanOut222;
wire [7:0] nOut13_15;
wire [7:0] nScanOut223;
wire [7:0] nOut14_0;
wire [7:0] nScanOut224;
wire [7:0] nOut14_1;
wire [7:0] nScanOut225;
wire [7:0] nOut14_2;
wire [7:0] nScanOut226;
wire [7:0] nOut14_3;
wire [7:0] nScanOut227;
wire [7:0] nOut14_4;
wire [7:0] nScanOut228;
wire [7:0] nOut14_5;
wire [7:0] nScanOut229;
wire [7:0] nOut14_6;
wire [7:0] nScanOut230;
wire [7:0] nOut14_7;
wire [7:0] nScanOut231;
wire [7:0] nOut14_8;
wire [7:0] nScanOut232;
wire [7:0] nOut14_9;
wire [7:0] nScanOut233;
wire [7:0] nOut14_10;
wire [7:0] nScanOut234;
wire [7:0] nOut14_11;
wire [7:0] nScanOut235;
wire [7:0] nOut14_12;
wire [7:0] nScanOut236;
wire [7:0] nOut14_13;
wire [7:0] nScanOut237;
wire [7:0] nOut14_14;
wire [7:0] nScanOut238;
wire [7:0] nOut14_15;
wire [7:0] nScanOut239;
wire [7:0] nOut15_0;
wire [7:0] nScanOut240;
wire [7:0] nOut15_1;
wire [7:0] nScanOut241;
wire [7:0] nOut15_2;
wire [7:0] nScanOut242;
wire [7:0] nOut15_3;
wire [7:0] nScanOut243;
wire [7:0] nOut15_4;
wire [7:0] nScanOut244;
wire [7:0] nOut15_5;
wire [7:0] nScanOut245;
wire [7:0] nOut15_6;
wire [7:0] nScanOut246;
wire [7:0] nOut15_7;
wire [7:0] nScanOut247;
wire [7:0] nOut15_8;
wire [7:0] nScanOut248;
wire [7:0] nOut15_9;
wire [7:0] nScanOut249;
wire [7:0] nOut15_10;
wire [7:0] nScanOut250;
wire [7:0] nOut15_11;
wire [7:0] nScanOut251;
wire [7:0] nOut15_12;
wire [7:0] nScanOut252;
wire [7:0] nOut15_13;
wire [7:0] nScanOut253;
wire [7:0] nOut15_14;
wire [7:0] nScanOut254;
wire [7:0] nOut15_15;
wire [7:0] nScanOut255;
wire [0:0] nEnable;
wire [0:0] nScanEnable;
wire [7:0] nScanOut256;
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_0), .ScanIn(nScanOut1), .ScanOut(nScanOut0), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_1), .ScanIn(nScanOut2), .ScanOut(nScanOut1), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_2), .ScanIn(nScanOut3), .ScanOut(nScanOut2), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_3), .ScanIn(nScanOut4), .ScanOut(nScanOut3), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_4), .ScanIn(nScanOut5), .ScanOut(nScanOut4), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_5), .ScanIn(nScanOut6), .ScanOut(nScanOut5), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_6), .ScanIn(nScanOut7), .ScanOut(nScanOut6), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_7), .ScanIn(nScanOut8), .ScanOut(nScanOut7), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_8), .ScanIn(nScanOut9), .ScanOut(nScanOut8), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_9), .ScanIn(nScanOut10), .ScanOut(nScanOut9), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_10), .ScanIn(nScanOut11), .ScanOut(nScanOut10), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_11), .ScanIn(nScanOut12), .ScanOut(nScanOut11), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_12), .ScanIn(nScanOut13), .ScanOut(nScanOut12), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_13), .ScanIn(nScanOut14), .ScanOut(nScanOut13), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_14), .ScanIn(nScanOut15), .ScanOut(nScanOut14), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_15), .ScanIn(nScanOut16), .ScanOut(nScanOut15), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_0), .ScanIn(nScanOut17), .ScanOut(nScanOut16), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_1), .NorthIn(nOut1_0), .SouthIn(nOut1_2), .EastIn(nOut2_1), .WestIn(nOut0_1), .ScanIn(nScanOut18), .ScanOut(nScanOut17), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_2), .NorthIn(nOut1_1), .SouthIn(nOut1_3), .EastIn(nOut2_2), .WestIn(nOut0_2), .ScanIn(nScanOut19), .ScanOut(nScanOut18), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_3), .NorthIn(nOut1_2), .SouthIn(nOut1_4), .EastIn(nOut2_3), .WestIn(nOut0_3), .ScanIn(nScanOut20), .ScanOut(nScanOut19), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_4), .NorthIn(nOut1_3), .SouthIn(nOut1_5), .EastIn(nOut2_4), .WestIn(nOut0_4), .ScanIn(nScanOut21), .ScanOut(nScanOut20), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_5), .NorthIn(nOut1_4), .SouthIn(nOut1_6), .EastIn(nOut2_5), .WestIn(nOut0_5), .ScanIn(nScanOut22), .ScanOut(nScanOut21), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_6), .NorthIn(nOut1_5), .SouthIn(nOut1_7), .EastIn(nOut2_6), .WestIn(nOut0_6), .ScanIn(nScanOut23), .ScanOut(nScanOut22), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_7), .NorthIn(nOut1_6), .SouthIn(nOut1_8), .EastIn(nOut2_7), .WestIn(nOut0_7), .ScanIn(nScanOut24), .ScanOut(nScanOut23), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_8), .NorthIn(nOut1_7), .SouthIn(nOut1_9), .EastIn(nOut2_8), .WestIn(nOut0_8), .ScanIn(nScanOut25), .ScanOut(nScanOut24), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_9), .NorthIn(nOut1_8), .SouthIn(nOut1_10), .EastIn(nOut2_9), .WestIn(nOut0_9), .ScanIn(nScanOut26), .ScanOut(nScanOut25), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_10), .NorthIn(nOut1_9), .SouthIn(nOut1_11), .EastIn(nOut2_10), .WestIn(nOut0_10), .ScanIn(nScanOut27), .ScanOut(nScanOut26), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_11), .NorthIn(nOut1_10), .SouthIn(nOut1_12), .EastIn(nOut2_11), .WestIn(nOut0_11), .ScanIn(nScanOut28), .ScanOut(nScanOut27), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_12), .NorthIn(nOut1_11), .SouthIn(nOut1_13), .EastIn(nOut2_12), .WestIn(nOut0_12), .ScanIn(nScanOut29), .ScanOut(nScanOut28), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_13), .NorthIn(nOut1_12), .SouthIn(nOut1_14), .EastIn(nOut2_13), .WestIn(nOut0_13), .ScanIn(nScanOut30), .ScanOut(nScanOut29), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_14), .NorthIn(nOut1_13), .SouthIn(nOut1_15), .EastIn(nOut2_14), .WestIn(nOut0_14), .ScanIn(nScanOut31), .ScanOut(nScanOut30), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_15), .ScanIn(nScanOut32), .ScanOut(nScanOut31), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_0), .ScanIn(nScanOut33), .ScanOut(nScanOut32), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_1), .NorthIn(nOut2_0), .SouthIn(nOut2_2), .EastIn(nOut3_1), .WestIn(nOut1_1), .ScanIn(nScanOut34), .ScanOut(nScanOut33), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_2), .NorthIn(nOut2_1), .SouthIn(nOut2_3), .EastIn(nOut3_2), .WestIn(nOut1_2), .ScanIn(nScanOut35), .ScanOut(nScanOut34), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_3), .NorthIn(nOut2_2), .SouthIn(nOut2_4), .EastIn(nOut3_3), .WestIn(nOut1_3), .ScanIn(nScanOut36), .ScanOut(nScanOut35), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_4), .NorthIn(nOut2_3), .SouthIn(nOut2_5), .EastIn(nOut3_4), .WestIn(nOut1_4), .ScanIn(nScanOut37), .ScanOut(nScanOut36), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_5), .NorthIn(nOut2_4), .SouthIn(nOut2_6), .EastIn(nOut3_5), .WestIn(nOut1_5), .ScanIn(nScanOut38), .ScanOut(nScanOut37), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_6), .NorthIn(nOut2_5), .SouthIn(nOut2_7), .EastIn(nOut3_6), .WestIn(nOut1_6), .ScanIn(nScanOut39), .ScanOut(nScanOut38), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_7), .NorthIn(nOut2_6), .SouthIn(nOut2_8), .EastIn(nOut3_7), .WestIn(nOut1_7), .ScanIn(nScanOut40), .ScanOut(nScanOut39), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_8), .NorthIn(nOut2_7), .SouthIn(nOut2_9), .EastIn(nOut3_8), .WestIn(nOut1_8), .ScanIn(nScanOut41), .ScanOut(nScanOut40), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_9), .NorthIn(nOut2_8), .SouthIn(nOut2_10), .EastIn(nOut3_9), .WestIn(nOut1_9), .ScanIn(nScanOut42), .ScanOut(nScanOut41), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_10), .NorthIn(nOut2_9), .SouthIn(nOut2_11), .EastIn(nOut3_10), .WestIn(nOut1_10), .ScanIn(nScanOut43), .ScanOut(nScanOut42), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_11), .NorthIn(nOut2_10), .SouthIn(nOut2_12), .EastIn(nOut3_11), .WestIn(nOut1_11), .ScanIn(nScanOut44), .ScanOut(nScanOut43), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_12), .NorthIn(nOut2_11), .SouthIn(nOut2_13), .EastIn(nOut3_12), .WestIn(nOut1_12), .ScanIn(nScanOut45), .ScanOut(nScanOut44), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_13), .NorthIn(nOut2_12), .SouthIn(nOut2_14), .EastIn(nOut3_13), .WestIn(nOut1_13), .ScanIn(nScanOut46), .ScanOut(nScanOut45), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_14), .NorthIn(nOut2_13), .SouthIn(nOut2_15), .EastIn(nOut3_14), .WestIn(nOut1_14), .ScanIn(nScanOut47), .ScanOut(nScanOut46), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_15), .ScanIn(nScanOut48), .ScanOut(nScanOut47), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_0), .ScanIn(nScanOut49), .ScanOut(nScanOut48), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_1), .NorthIn(nOut3_0), .SouthIn(nOut3_2), .EastIn(nOut4_1), .WestIn(nOut2_1), .ScanIn(nScanOut50), .ScanOut(nScanOut49), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_2), .NorthIn(nOut3_1), .SouthIn(nOut3_3), .EastIn(nOut4_2), .WestIn(nOut2_2), .ScanIn(nScanOut51), .ScanOut(nScanOut50), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_3), .NorthIn(nOut3_2), .SouthIn(nOut3_4), .EastIn(nOut4_3), .WestIn(nOut2_3), .ScanIn(nScanOut52), .ScanOut(nScanOut51), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_4), .NorthIn(nOut3_3), .SouthIn(nOut3_5), .EastIn(nOut4_4), .WestIn(nOut2_4), .ScanIn(nScanOut53), .ScanOut(nScanOut52), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_5), .NorthIn(nOut3_4), .SouthIn(nOut3_6), .EastIn(nOut4_5), .WestIn(nOut2_5), .ScanIn(nScanOut54), .ScanOut(nScanOut53), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_6), .NorthIn(nOut3_5), .SouthIn(nOut3_7), .EastIn(nOut4_6), .WestIn(nOut2_6), .ScanIn(nScanOut55), .ScanOut(nScanOut54), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_7), .NorthIn(nOut3_6), .SouthIn(nOut3_8), .EastIn(nOut4_7), .WestIn(nOut2_7), .ScanIn(nScanOut56), .ScanOut(nScanOut55), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_8), .NorthIn(nOut3_7), .SouthIn(nOut3_9), .EastIn(nOut4_8), .WestIn(nOut2_8), .ScanIn(nScanOut57), .ScanOut(nScanOut56), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_9), .NorthIn(nOut3_8), .SouthIn(nOut3_10), .EastIn(nOut4_9), .WestIn(nOut2_9), .ScanIn(nScanOut58), .ScanOut(nScanOut57), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_10), .NorthIn(nOut3_9), .SouthIn(nOut3_11), .EastIn(nOut4_10), .WestIn(nOut2_10), .ScanIn(nScanOut59), .ScanOut(nScanOut58), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_11), .NorthIn(nOut3_10), .SouthIn(nOut3_12), .EastIn(nOut4_11), .WestIn(nOut2_11), .ScanIn(nScanOut60), .ScanOut(nScanOut59), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_12), .NorthIn(nOut3_11), .SouthIn(nOut3_13), .EastIn(nOut4_12), .WestIn(nOut2_12), .ScanIn(nScanOut61), .ScanOut(nScanOut60), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_13), .NorthIn(nOut3_12), .SouthIn(nOut3_14), .EastIn(nOut4_13), .WestIn(nOut2_13), .ScanIn(nScanOut62), .ScanOut(nScanOut61), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_14), .NorthIn(nOut3_13), .SouthIn(nOut3_15), .EastIn(nOut4_14), .WestIn(nOut2_14), .ScanIn(nScanOut63), .ScanOut(nScanOut62), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_15), .ScanIn(nScanOut64), .ScanOut(nScanOut63), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_64 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_0), .ScanIn(nScanOut65), .ScanOut(nScanOut64), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_65 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_1), .NorthIn(nOut4_0), .SouthIn(nOut4_2), .EastIn(nOut5_1), .WestIn(nOut3_1), .ScanIn(nScanOut66), .ScanOut(nScanOut65), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_66 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_2), .NorthIn(nOut4_1), .SouthIn(nOut4_3), .EastIn(nOut5_2), .WestIn(nOut3_2), .ScanIn(nScanOut67), .ScanOut(nScanOut66), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_67 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_3), .NorthIn(nOut4_2), .SouthIn(nOut4_4), .EastIn(nOut5_3), .WestIn(nOut3_3), .ScanIn(nScanOut68), .ScanOut(nScanOut67), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_68 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_4), .NorthIn(nOut4_3), .SouthIn(nOut4_5), .EastIn(nOut5_4), .WestIn(nOut3_4), .ScanIn(nScanOut69), .ScanOut(nScanOut68), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_69 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_5), .NorthIn(nOut4_4), .SouthIn(nOut4_6), .EastIn(nOut5_5), .WestIn(nOut3_5), .ScanIn(nScanOut70), .ScanOut(nScanOut69), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_70 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_6), .NorthIn(nOut4_5), .SouthIn(nOut4_7), .EastIn(nOut5_6), .WestIn(nOut3_6), .ScanIn(nScanOut71), .ScanOut(nScanOut70), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_71 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_7), .NorthIn(nOut4_6), .SouthIn(nOut4_8), .EastIn(nOut5_7), .WestIn(nOut3_7), .ScanIn(nScanOut72), .ScanOut(nScanOut71), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_72 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_8), .NorthIn(nOut4_7), .SouthIn(nOut4_9), .EastIn(nOut5_8), .WestIn(nOut3_8), .ScanIn(nScanOut73), .ScanOut(nScanOut72), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_73 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_9), .NorthIn(nOut4_8), .SouthIn(nOut4_10), .EastIn(nOut5_9), .WestIn(nOut3_9), .ScanIn(nScanOut74), .ScanOut(nScanOut73), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_74 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_10), .NorthIn(nOut4_9), .SouthIn(nOut4_11), .EastIn(nOut5_10), .WestIn(nOut3_10), .ScanIn(nScanOut75), .ScanOut(nScanOut74), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_75 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_11), .NorthIn(nOut4_10), .SouthIn(nOut4_12), .EastIn(nOut5_11), .WestIn(nOut3_11), .ScanIn(nScanOut76), .ScanOut(nScanOut75), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_76 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_12), .NorthIn(nOut4_11), .SouthIn(nOut4_13), .EastIn(nOut5_12), .WestIn(nOut3_12), .ScanIn(nScanOut77), .ScanOut(nScanOut76), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_77 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_13), .NorthIn(nOut4_12), .SouthIn(nOut4_14), .EastIn(nOut5_13), .WestIn(nOut3_13), .ScanIn(nScanOut78), .ScanOut(nScanOut77), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_78 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_14), .NorthIn(nOut4_13), .SouthIn(nOut4_15), .EastIn(nOut5_14), .WestIn(nOut3_14), .ScanIn(nScanOut79), .ScanOut(nScanOut78), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_79 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_15), .ScanIn(nScanOut80), .ScanOut(nScanOut79), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_80 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_0), .ScanIn(nScanOut81), .ScanOut(nScanOut80), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_81 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_1), .NorthIn(nOut5_0), .SouthIn(nOut5_2), .EastIn(nOut6_1), .WestIn(nOut4_1), .ScanIn(nScanOut82), .ScanOut(nScanOut81), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_82 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_2), .NorthIn(nOut5_1), .SouthIn(nOut5_3), .EastIn(nOut6_2), .WestIn(nOut4_2), .ScanIn(nScanOut83), .ScanOut(nScanOut82), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_83 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_3), .NorthIn(nOut5_2), .SouthIn(nOut5_4), .EastIn(nOut6_3), .WestIn(nOut4_3), .ScanIn(nScanOut84), .ScanOut(nScanOut83), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_84 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_4), .NorthIn(nOut5_3), .SouthIn(nOut5_5), .EastIn(nOut6_4), .WestIn(nOut4_4), .ScanIn(nScanOut85), .ScanOut(nScanOut84), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_85 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_5), .NorthIn(nOut5_4), .SouthIn(nOut5_6), .EastIn(nOut6_5), .WestIn(nOut4_5), .ScanIn(nScanOut86), .ScanOut(nScanOut85), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_86 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_6), .NorthIn(nOut5_5), .SouthIn(nOut5_7), .EastIn(nOut6_6), .WestIn(nOut4_6), .ScanIn(nScanOut87), .ScanOut(nScanOut86), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_87 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_7), .NorthIn(nOut5_6), .SouthIn(nOut5_8), .EastIn(nOut6_7), .WestIn(nOut4_7), .ScanIn(nScanOut88), .ScanOut(nScanOut87), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_88 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_8), .NorthIn(nOut5_7), .SouthIn(nOut5_9), .EastIn(nOut6_8), .WestIn(nOut4_8), .ScanIn(nScanOut89), .ScanOut(nScanOut88), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_89 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_9), .NorthIn(nOut5_8), .SouthIn(nOut5_10), .EastIn(nOut6_9), .WestIn(nOut4_9), .ScanIn(nScanOut90), .ScanOut(nScanOut89), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_90 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_10), .NorthIn(nOut5_9), .SouthIn(nOut5_11), .EastIn(nOut6_10), .WestIn(nOut4_10), .ScanIn(nScanOut91), .ScanOut(nScanOut90), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_91 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_11), .NorthIn(nOut5_10), .SouthIn(nOut5_12), .EastIn(nOut6_11), .WestIn(nOut4_11), .ScanIn(nScanOut92), .ScanOut(nScanOut91), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_92 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_12), .NorthIn(nOut5_11), .SouthIn(nOut5_13), .EastIn(nOut6_12), .WestIn(nOut4_12), .ScanIn(nScanOut93), .ScanOut(nScanOut92), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_93 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_13), .NorthIn(nOut5_12), .SouthIn(nOut5_14), .EastIn(nOut6_13), .WestIn(nOut4_13), .ScanIn(nScanOut94), .ScanOut(nScanOut93), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_94 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_14), .NorthIn(nOut5_13), .SouthIn(nOut5_15), .EastIn(nOut6_14), .WestIn(nOut4_14), .ScanIn(nScanOut95), .ScanOut(nScanOut94), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_95 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_15), .ScanIn(nScanOut96), .ScanOut(nScanOut95), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_96 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_0), .ScanIn(nScanOut97), .ScanOut(nScanOut96), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_97 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_1), .NorthIn(nOut6_0), .SouthIn(nOut6_2), .EastIn(nOut7_1), .WestIn(nOut5_1), .ScanIn(nScanOut98), .ScanOut(nScanOut97), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_98 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_2), .NorthIn(nOut6_1), .SouthIn(nOut6_3), .EastIn(nOut7_2), .WestIn(nOut5_2), .ScanIn(nScanOut99), .ScanOut(nScanOut98), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_99 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_3), .NorthIn(nOut6_2), .SouthIn(nOut6_4), .EastIn(nOut7_3), .WestIn(nOut5_3), .ScanIn(nScanOut100), .ScanOut(nScanOut99), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_100 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_4), .NorthIn(nOut6_3), .SouthIn(nOut6_5), .EastIn(nOut7_4), .WestIn(nOut5_4), .ScanIn(nScanOut101), .ScanOut(nScanOut100), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_101 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_5), .NorthIn(nOut6_4), .SouthIn(nOut6_6), .EastIn(nOut7_5), .WestIn(nOut5_5), .ScanIn(nScanOut102), .ScanOut(nScanOut101), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_102 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_6), .NorthIn(nOut6_5), .SouthIn(nOut6_7), .EastIn(nOut7_6), .WestIn(nOut5_6), .ScanIn(nScanOut103), .ScanOut(nScanOut102), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_103 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_7), .NorthIn(nOut6_6), .SouthIn(nOut6_8), .EastIn(nOut7_7), .WestIn(nOut5_7), .ScanIn(nScanOut104), .ScanOut(nScanOut103), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_104 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_8), .NorthIn(nOut6_7), .SouthIn(nOut6_9), .EastIn(nOut7_8), .WestIn(nOut5_8), .ScanIn(nScanOut105), .ScanOut(nScanOut104), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_105 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_9), .NorthIn(nOut6_8), .SouthIn(nOut6_10), .EastIn(nOut7_9), .WestIn(nOut5_9), .ScanIn(nScanOut106), .ScanOut(nScanOut105), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_106 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_10), .NorthIn(nOut6_9), .SouthIn(nOut6_11), .EastIn(nOut7_10), .WestIn(nOut5_10), .ScanIn(nScanOut107), .ScanOut(nScanOut106), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_107 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_11), .NorthIn(nOut6_10), .SouthIn(nOut6_12), .EastIn(nOut7_11), .WestIn(nOut5_11), .ScanIn(nScanOut108), .ScanOut(nScanOut107), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_108 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_12), .NorthIn(nOut6_11), .SouthIn(nOut6_13), .EastIn(nOut7_12), .WestIn(nOut5_12), .ScanIn(nScanOut109), .ScanOut(nScanOut108), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_109 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_13), .NorthIn(nOut6_12), .SouthIn(nOut6_14), .EastIn(nOut7_13), .WestIn(nOut5_13), .ScanIn(nScanOut110), .ScanOut(nScanOut109), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_110 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_14), .NorthIn(nOut6_13), .SouthIn(nOut6_15), .EastIn(nOut7_14), .WestIn(nOut5_14), .ScanIn(nScanOut111), .ScanOut(nScanOut110), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_111 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_15), .ScanIn(nScanOut112), .ScanOut(nScanOut111), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_112 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_0), .ScanIn(nScanOut113), .ScanOut(nScanOut112), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_113 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_1), .NorthIn(nOut7_0), .SouthIn(nOut7_2), .EastIn(nOut8_1), .WestIn(nOut6_1), .ScanIn(nScanOut114), .ScanOut(nScanOut113), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_114 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_2), .NorthIn(nOut7_1), .SouthIn(nOut7_3), .EastIn(nOut8_2), .WestIn(nOut6_2), .ScanIn(nScanOut115), .ScanOut(nScanOut114), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_115 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_3), .NorthIn(nOut7_2), .SouthIn(nOut7_4), .EastIn(nOut8_3), .WestIn(nOut6_3), .ScanIn(nScanOut116), .ScanOut(nScanOut115), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_116 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_4), .NorthIn(nOut7_3), .SouthIn(nOut7_5), .EastIn(nOut8_4), .WestIn(nOut6_4), .ScanIn(nScanOut117), .ScanOut(nScanOut116), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_117 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_5), .NorthIn(nOut7_4), .SouthIn(nOut7_6), .EastIn(nOut8_5), .WestIn(nOut6_5), .ScanIn(nScanOut118), .ScanOut(nScanOut117), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_118 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_6), .NorthIn(nOut7_5), .SouthIn(nOut7_7), .EastIn(nOut8_6), .WestIn(nOut6_6), .ScanIn(nScanOut119), .ScanOut(nScanOut118), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_119 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_7), .NorthIn(nOut7_6), .SouthIn(nOut7_8), .EastIn(nOut8_7), .WestIn(nOut6_7), .ScanIn(nScanOut120), .ScanOut(nScanOut119), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_120 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_8), .NorthIn(nOut7_7), .SouthIn(nOut7_9), .EastIn(nOut8_8), .WestIn(nOut6_8), .ScanIn(nScanOut121), .ScanOut(nScanOut120), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_121 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_9), .NorthIn(nOut7_8), .SouthIn(nOut7_10), .EastIn(nOut8_9), .WestIn(nOut6_9), .ScanIn(nScanOut122), .ScanOut(nScanOut121), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_122 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_10), .NorthIn(nOut7_9), .SouthIn(nOut7_11), .EastIn(nOut8_10), .WestIn(nOut6_10), .ScanIn(nScanOut123), .ScanOut(nScanOut122), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_123 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_11), .NorthIn(nOut7_10), .SouthIn(nOut7_12), .EastIn(nOut8_11), .WestIn(nOut6_11), .ScanIn(nScanOut124), .ScanOut(nScanOut123), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_124 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_12), .NorthIn(nOut7_11), .SouthIn(nOut7_13), .EastIn(nOut8_12), .WestIn(nOut6_12), .ScanIn(nScanOut125), .ScanOut(nScanOut124), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_125 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_13), .NorthIn(nOut7_12), .SouthIn(nOut7_14), .EastIn(nOut8_13), .WestIn(nOut6_13), .ScanIn(nScanOut126), .ScanOut(nScanOut125), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_126 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut7_14), .NorthIn(nOut7_13), .SouthIn(nOut7_15), .EastIn(nOut8_14), .WestIn(nOut6_14), .ScanIn(nScanOut127), .ScanOut(nScanOut126), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_127 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_15), .ScanIn(nScanOut128), .ScanOut(nScanOut127), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_128 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut8_0), .ScanIn(nScanOut129), .ScanOut(nScanOut128), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_129 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_1), .NorthIn(nOut8_0), .SouthIn(nOut8_2), .EastIn(nOut9_1), .WestIn(nOut7_1), .ScanIn(nScanOut130), .ScanOut(nScanOut129), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_130 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_2), .NorthIn(nOut8_1), .SouthIn(nOut8_3), .EastIn(nOut9_2), .WestIn(nOut7_2), .ScanIn(nScanOut131), .ScanOut(nScanOut130), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_131 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_3), .NorthIn(nOut8_2), .SouthIn(nOut8_4), .EastIn(nOut9_3), .WestIn(nOut7_3), .ScanIn(nScanOut132), .ScanOut(nScanOut131), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_132 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_4), .NorthIn(nOut8_3), .SouthIn(nOut8_5), .EastIn(nOut9_4), .WestIn(nOut7_4), .ScanIn(nScanOut133), .ScanOut(nScanOut132), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_133 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_5), .NorthIn(nOut8_4), .SouthIn(nOut8_6), .EastIn(nOut9_5), .WestIn(nOut7_5), .ScanIn(nScanOut134), .ScanOut(nScanOut133), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_134 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_6), .NorthIn(nOut8_5), .SouthIn(nOut8_7), .EastIn(nOut9_6), .WestIn(nOut7_6), .ScanIn(nScanOut135), .ScanOut(nScanOut134), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_135 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_7), .NorthIn(nOut8_6), .SouthIn(nOut8_8), .EastIn(nOut9_7), .WestIn(nOut7_7), .ScanIn(nScanOut136), .ScanOut(nScanOut135), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_136 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_8), .NorthIn(nOut8_7), .SouthIn(nOut8_9), .EastIn(nOut9_8), .WestIn(nOut7_8), .ScanIn(nScanOut137), .ScanOut(nScanOut136), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_137 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_9), .NorthIn(nOut8_8), .SouthIn(nOut8_10), .EastIn(nOut9_9), .WestIn(nOut7_9), .ScanIn(nScanOut138), .ScanOut(nScanOut137), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_138 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_10), .NorthIn(nOut8_9), .SouthIn(nOut8_11), .EastIn(nOut9_10), .WestIn(nOut7_10), .ScanIn(nScanOut139), .ScanOut(nScanOut138), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_139 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_11), .NorthIn(nOut8_10), .SouthIn(nOut8_12), .EastIn(nOut9_11), .WestIn(nOut7_11), .ScanIn(nScanOut140), .ScanOut(nScanOut139), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_140 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_12), .NorthIn(nOut8_11), .SouthIn(nOut8_13), .EastIn(nOut9_12), .WestIn(nOut7_12), .ScanIn(nScanOut141), .ScanOut(nScanOut140), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_141 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_13), .NorthIn(nOut8_12), .SouthIn(nOut8_14), .EastIn(nOut9_13), .WestIn(nOut7_13), .ScanIn(nScanOut142), .ScanOut(nScanOut141), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_142 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut8_14), .NorthIn(nOut8_13), .SouthIn(nOut8_15), .EastIn(nOut9_14), .WestIn(nOut7_14), .ScanIn(nScanOut143), .ScanOut(nScanOut142), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_143 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut8_15), .ScanIn(nScanOut144), .ScanOut(nScanOut143), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_144 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut9_0), .ScanIn(nScanOut145), .ScanOut(nScanOut144), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_145 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_1), .NorthIn(nOut9_0), .SouthIn(nOut9_2), .EastIn(nOut10_1), .WestIn(nOut8_1), .ScanIn(nScanOut146), .ScanOut(nScanOut145), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_146 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_2), .NorthIn(nOut9_1), .SouthIn(nOut9_3), .EastIn(nOut10_2), .WestIn(nOut8_2), .ScanIn(nScanOut147), .ScanOut(nScanOut146), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_147 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_3), .NorthIn(nOut9_2), .SouthIn(nOut9_4), .EastIn(nOut10_3), .WestIn(nOut8_3), .ScanIn(nScanOut148), .ScanOut(nScanOut147), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_148 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_4), .NorthIn(nOut9_3), .SouthIn(nOut9_5), .EastIn(nOut10_4), .WestIn(nOut8_4), .ScanIn(nScanOut149), .ScanOut(nScanOut148), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_149 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_5), .NorthIn(nOut9_4), .SouthIn(nOut9_6), .EastIn(nOut10_5), .WestIn(nOut8_5), .ScanIn(nScanOut150), .ScanOut(nScanOut149), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_150 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_6), .NorthIn(nOut9_5), .SouthIn(nOut9_7), .EastIn(nOut10_6), .WestIn(nOut8_6), .ScanIn(nScanOut151), .ScanOut(nScanOut150), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_151 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_7), .NorthIn(nOut9_6), .SouthIn(nOut9_8), .EastIn(nOut10_7), .WestIn(nOut8_7), .ScanIn(nScanOut152), .ScanOut(nScanOut151), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_152 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_8), .NorthIn(nOut9_7), .SouthIn(nOut9_9), .EastIn(nOut10_8), .WestIn(nOut8_8), .ScanIn(nScanOut153), .ScanOut(nScanOut152), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_153 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_9), .NorthIn(nOut9_8), .SouthIn(nOut9_10), .EastIn(nOut10_9), .WestIn(nOut8_9), .ScanIn(nScanOut154), .ScanOut(nScanOut153), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_154 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_10), .NorthIn(nOut9_9), .SouthIn(nOut9_11), .EastIn(nOut10_10), .WestIn(nOut8_10), .ScanIn(nScanOut155), .ScanOut(nScanOut154), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_155 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_11), .NorthIn(nOut9_10), .SouthIn(nOut9_12), .EastIn(nOut10_11), .WestIn(nOut8_11), .ScanIn(nScanOut156), .ScanOut(nScanOut155), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_156 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_12), .NorthIn(nOut9_11), .SouthIn(nOut9_13), .EastIn(nOut10_12), .WestIn(nOut8_12), .ScanIn(nScanOut157), .ScanOut(nScanOut156), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_157 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_13), .NorthIn(nOut9_12), .SouthIn(nOut9_14), .EastIn(nOut10_13), .WestIn(nOut8_13), .ScanIn(nScanOut158), .ScanOut(nScanOut157), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_158 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut9_14), .NorthIn(nOut9_13), .SouthIn(nOut9_15), .EastIn(nOut10_14), .WestIn(nOut8_14), .ScanIn(nScanOut159), .ScanOut(nScanOut158), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_159 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut9_15), .ScanIn(nScanOut160), .ScanOut(nScanOut159), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_160 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut10_0), .ScanIn(nScanOut161), .ScanOut(nScanOut160), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_161 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_1), .NorthIn(nOut10_0), .SouthIn(nOut10_2), .EastIn(nOut11_1), .WestIn(nOut9_1), .ScanIn(nScanOut162), .ScanOut(nScanOut161), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_162 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_2), .NorthIn(nOut10_1), .SouthIn(nOut10_3), .EastIn(nOut11_2), .WestIn(nOut9_2), .ScanIn(nScanOut163), .ScanOut(nScanOut162), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_163 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_3), .NorthIn(nOut10_2), .SouthIn(nOut10_4), .EastIn(nOut11_3), .WestIn(nOut9_3), .ScanIn(nScanOut164), .ScanOut(nScanOut163), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_164 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_4), .NorthIn(nOut10_3), .SouthIn(nOut10_5), .EastIn(nOut11_4), .WestIn(nOut9_4), .ScanIn(nScanOut165), .ScanOut(nScanOut164), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_165 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_5), .NorthIn(nOut10_4), .SouthIn(nOut10_6), .EastIn(nOut11_5), .WestIn(nOut9_5), .ScanIn(nScanOut166), .ScanOut(nScanOut165), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_166 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_6), .NorthIn(nOut10_5), .SouthIn(nOut10_7), .EastIn(nOut11_6), .WestIn(nOut9_6), .ScanIn(nScanOut167), .ScanOut(nScanOut166), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_167 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_7), .NorthIn(nOut10_6), .SouthIn(nOut10_8), .EastIn(nOut11_7), .WestIn(nOut9_7), .ScanIn(nScanOut168), .ScanOut(nScanOut167), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_168 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_8), .NorthIn(nOut10_7), .SouthIn(nOut10_9), .EastIn(nOut11_8), .WestIn(nOut9_8), .ScanIn(nScanOut169), .ScanOut(nScanOut168), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_169 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_9), .NorthIn(nOut10_8), .SouthIn(nOut10_10), .EastIn(nOut11_9), .WestIn(nOut9_9), .ScanIn(nScanOut170), .ScanOut(nScanOut169), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_170 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_10), .NorthIn(nOut10_9), .SouthIn(nOut10_11), .EastIn(nOut11_10), .WestIn(nOut9_10), .ScanIn(nScanOut171), .ScanOut(nScanOut170), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_171 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_11), .NorthIn(nOut10_10), .SouthIn(nOut10_12), .EastIn(nOut11_11), .WestIn(nOut9_11), .ScanIn(nScanOut172), .ScanOut(nScanOut171), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_172 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_12), .NorthIn(nOut10_11), .SouthIn(nOut10_13), .EastIn(nOut11_12), .WestIn(nOut9_12), .ScanIn(nScanOut173), .ScanOut(nScanOut172), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_173 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_13), .NorthIn(nOut10_12), .SouthIn(nOut10_14), .EastIn(nOut11_13), .WestIn(nOut9_13), .ScanIn(nScanOut174), .ScanOut(nScanOut173), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_174 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut10_14), .NorthIn(nOut10_13), .SouthIn(nOut10_15), .EastIn(nOut11_14), .WestIn(nOut9_14), .ScanIn(nScanOut175), .ScanOut(nScanOut174), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_175 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut10_15), .ScanIn(nScanOut176), .ScanOut(nScanOut175), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_176 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut11_0), .ScanIn(nScanOut177), .ScanOut(nScanOut176), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_177 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_1), .NorthIn(nOut11_0), .SouthIn(nOut11_2), .EastIn(nOut12_1), .WestIn(nOut10_1), .ScanIn(nScanOut178), .ScanOut(nScanOut177), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_178 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_2), .NorthIn(nOut11_1), .SouthIn(nOut11_3), .EastIn(nOut12_2), .WestIn(nOut10_2), .ScanIn(nScanOut179), .ScanOut(nScanOut178), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_179 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_3), .NorthIn(nOut11_2), .SouthIn(nOut11_4), .EastIn(nOut12_3), .WestIn(nOut10_3), .ScanIn(nScanOut180), .ScanOut(nScanOut179), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_180 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_4), .NorthIn(nOut11_3), .SouthIn(nOut11_5), .EastIn(nOut12_4), .WestIn(nOut10_4), .ScanIn(nScanOut181), .ScanOut(nScanOut180), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_181 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_5), .NorthIn(nOut11_4), .SouthIn(nOut11_6), .EastIn(nOut12_5), .WestIn(nOut10_5), .ScanIn(nScanOut182), .ScanOut(nScanOut181), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_182 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_6), .NorthIn(nOut11_5), .SouthIn(nOut11_7), .EastIn(nOut12_6), .WestIn(nOut10_6), .ScanIn(nScanOut183), .ScanOut(nScanOut182), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_183 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_7), .NorthIn(nOut11_6), .SouthIn(nOut11_8), .EastIn(nOut12_7), .WestIn(nOut10_7), .ScanIn(nScanOut184), .ScanOut(nScanOut183), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_184 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_8), .NorthIn(nOut11_7), .SouthIn(nOut11_9), .EastIn(nOut12_8), .WestIn(nOut10_8), .ScanIn(nScanOut185), .ScanOut(nScanOut184), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_185 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_9), .NorthIn(nOut11_8), .SouthIn(nOut11_10), .EastIn(nOut12_9), .WestIn(nOut10_9), .ScanIn(nScanOut186), .ScanOut(nScanOut185), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_186 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_10), .NorthIn(nOut11_9), .SouthIn(nOut11_11), .EastIn(nOut12_10), .WestIn(nOut10_10), .ScanIn(nScanOut187), .ScanOut(nScanOut186), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_187 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_11), .NorthIn(nOut11_10), .SouthIn(nOut11_12), .EastIn(nOut12_11), .WestIn(nOut10_11), .ScanIn(nScanOut188), .ScanOut(nScanOut187), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_188 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_12), .NorthIn(nOut11_11), .SouthIn(nOut11_13), .EastIn(nOut12_12), .WestIn(nOut10_12), .ScanIn(nScanOut189), .ScanOut(nScanOut188), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_189 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_13), .NorthIn(nOut11_12), .SouthIn(nOut11_14), .EastIn(nOut12_13), .WestIn(nOut10_13), .ScanIn(nScanOut190), .ScanOut(nScanOut189), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_190 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut11_14), .NorthIn(nOut11_13), .SouthIn(nOut11_15), .EastIn(nOut12_14), .WestIn(nOut10_14), .ScanIn(nScanOut191), .ScanOut(nScanOut190), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_191 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut11_15), .ScanIn(nScanOut192), .ScanOut(nScanOut191), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_192 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut12_0), .ScanIn(nScanOut193), .ScanOut(nScanOut192), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_193 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_1), .NorthIn(nOut12_0), .SouthIn(nOut12_2), .EastIn(nOut13_1), .WestIn(nOut11_1), .ScanIn(nScanOut194), .ScanOut(nScanOut193), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_194 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_2), .NorthIn(nOut12_1), .SouthIn(nOut12_3), .EastIn(nOut13_2), .WestIn(nOut11_2), .ScanIn(nScanOut195), .ScanOut(nScanOut194), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_195 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_3), .NorthIn(nOut12_2), .SouthIn(nOut12_4), .EastIn(nOut13_3), .WestIn(nOut11_3), .ScanIn(nScanOut196), .ScanOut(nScanOut195), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_196 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_4), .NorthIn(nOut12_3), .SouthIn(nOut12_5), .EastIn(nOut13_4), .WestIn(nOut11_4), .ScanIn(nScanOut197), .ScanOut(nScanOut196), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_197 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_5), .NorthIn(nOut12_4), .SouthIn(nOut12_6), .EastIn(nOut13_5), .WestIn(nOut11_5), .ScanIn(nScanOut198), .ScanOut(nScanOut197), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_198 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_6), .NorthIn(nOut12_5), .SouthIn(nOut12_7), .EastIn(nOut13_6), .WestIn(nOut11_6), .ScanIn(nScanOut199), .ScanOut(nScanOut198), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_199 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_7), .NorthIn(nOut12_6), .SouthIn(nOut12_8), .EastIn(nOut13_7), .WestIn(nOut11_7), .ScanIn(nScanOut200), .ScanOut(nScanOut199), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_200 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_8), .NorthIn(nOut12_7), .SouthIn(nOut12_9), .EastIn(nOut13_8), .WestIn(nOut11_8), .ScanIn(nScanOut201), .ScanOut(nScanOut200), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_201 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_9), .NorthIn(nOut12_8), .SouthIn(nOut12_10), .EastIn(nOut13_9), .WestIn(nOut11_9), .ScanIn(nScanOut202), .ScanOut(nScanOut201), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_202 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_10), .NorthIn(nOut12_9), .SouthIn(nOut12_11), .EastIn(nOut13_10), .WestIn(nOut11_10), .ScanIn(nScanOut203), .ScanOut(nScanOut202), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_203 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_11), .NorthIn(nOut12_10), .SouthIn(nOut12_12), .EastIn(nOut13_11), .WestIn(nOut11_11), .ScanIn(nScanOut204), .ScanOut(nScanOut203), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_204 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_12), .NorthIn(nOut12_11), .SouthIn(nOut12_13), .EastIn(nOut13_12), .WestIn(nOut11_12), .ScanIn(nScanOut205), .ScanOut(nScanOut204), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_205 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_13), .NorthIn(nOut12_12), .SouthIn(nOut12_14), .EastIn(nOut13_13), .WestIn(nOut11_13), .ScanIn(nScanOut206), .ScanOut(nScanOut205), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_206 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut12_14), .NorthIn(nOut12_13), .SouthIn(nOut12_15), .EastIn(nOut13_14), .WestIn(nOut11_14), .ScanIn(nScanOut207), .ScanOut(nScanOut206), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_207 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut12_15), .ScanIn(nScanOut208), .ScanOut(nScanOut207), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_208 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut13_0), .ScanIn(nScanOut209), .ScanOut(nScanOut208), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_209 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_1), .NorthIn(nOut13_0), .SouthIn(nOut13_2), .EastIn(nOut14_1), .WestIn(nOut12_1), .ScanIn(nScanOut210), .ScanOut(nScanOut209), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_210 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_2), .NorthIn(nOut13_1), .SouthIn(nOut13_3), .EastIn(nOut14_2), .WestIn(nOut12_2), .ScanIn(nScanOut211), .ScanOut(nScanOut210), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_211 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_3), .NorthIn(nOut13_2), .SouthIn(nOut13_4), .EastIn(nOut14_3), .WestIn(nOut12_3), .ScanIn(nScanOut212), .ScanOut(nScanOut211), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_212 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_4), .NorthIn(nOut13_3), .SouthIn(nOut13_5), .EastIn(nOut14_4), .WestIn(nOut12_4), .ScanIn(nScanOut213), .ScanOut(nScanOut212), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_213 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_5), .NorthIn(nOut13_4), .SouthIn(nOut13_6), .EastIn(nOut14_5), .WestIn(nOut12_5), .ScanIn(nScanOut214), .ScanOut(nScanOut213), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_214 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_6), .NorthIn(nOut13_5), .SouthIn(nOut13_7), .EastIn(nOut14_6), .WestIn(nOut12_6), .ScanIn(nScanOut215), .ScanOut(nScanOut214), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_215 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_7), .NorthIn(nOut13_6), .SouthIn(nOut13_8), .EastIn(nOut14_7), .WestIn(nOut12_7), .ScanIn(nScanOut216), .ScanOut(nScanOut215), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_216 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_8), .NorthIn(nOut13_7), .SouthIn(nOut13_9), .EastIn(nOut14_8), .WestIn(nOut12_8), .ScanIn(nScanOut217), .ScanOut(nScanOut216), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_217 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_9), .NorthIn(nOut13_8), .SouthIn(nOut13_10), .EastIn(nOut14_9), .WestIn(nOut12_9), .ScanIn(nScanOut218), .ScanOut(nScanOut217), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_218 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_10), .NorthIn(nOut13_9), .SouthIn(nOut13_11), .EastIn(nOut14_10), .WestIn(nOut12_10), .ScanIn(nScanOut219), .ScanOut(nScanOut218), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_219 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_11), .NorthIn(nOut13_10), .SouthIn(nOut13_12), .EastIn(nOut14_11), .WestIn(nOut12_11), .ScanIn(nScanOut220), .ScanOut(nScanOut219), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_220 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_12), .NorthIn(nOut13_11), .SouthIn(nOut13_13), .EastIn(nOut14_12), .WestIn(nOut12_12), .ScanIn(nScanOut221), .ScanOut(nScanOut220), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_221 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_13), .NorthIn(nOut13_12), .SouthIn(nOut13_14), .EastIn(nOut14_13), .WestIn(nOut12_13), .ScanIn(nScanOut222), .ScanOut(nScanOut221), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_222 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut13_14), .NorthIn(nOut13_13), .SouthIn(nOut13_15), .EastIn(nOut14_14), .WestIn(nOut12_14), .ScanIn(nScanOut223), .ScanOut(nScanOut222), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_223 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut13_15), .ScanIn(nScanOut224), .ScanOut(nScanOut223), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_224 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut14_0), .ScanIn(nScanOut225), .ScanOut(nScanOut224), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_225 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_1), .NorthIn(nOut14_0), .SouthIn(nOut14_2), .EastIn(nOut15_1), .WestIn(nOut13_1), .ScanIn(nScanOut226), .ScanOut(nScanOut225), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_226 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_2), .NorthIn(nOut14_1), .SouthIn(nOut14_3), .EastIn(nOut15_2), .WestIn(nOut13_2), .ScanIn(nScanOut227), .ScanOut(nScanOut226), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_227 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_3), .NorthIn(nOut14_2), .SouthIn(nOut14_4), .EastIn(nOut15_3), .WestIn(nOut13_3), .ScanIn(nScanOut228), .ScanOut(nScanOut227), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_228 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_4), .NorthIn(nOut14_3), .SouthIn(nOut14_5), .EastIn(nOut15_4), .WestIn(nOut13_4), .ScanIn(nScanOut229), .ScanOut(nScanOut228), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_229 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_5), .NorthIn(nOut14_4), .SouthIn(nOut14_6), .EastIn(nOut15_5), .WestIn(nOut13_5), .ScanIn(nScanOut230), .ScanOut(nScanOut229), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_230 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_6), .NorthIn(nOut14_5), .SouthIn(nOut14_7), .EastIn(nOut15_6), .WestIn(nOut13_6), .ScanIn(nScanOut231), .ScanOut(nScanOut230), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_231 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_7), .NorthIn(nOut14_6), .SouthIn(nOut14_8), .EastIn(nOut15_7), .WestIn(nOut13_7), .ScanIn(nScanOut232), .ScanOut(nScanOut231), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_232 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_8), .NorthIn(nOut14_7), .SouthIn(nOut14_9), .EastIn(nOut15_8), .WestIn(nOut13_8), .ScanIn(nScanOut233), .ScanOut(nScanOut232), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_233 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_9), .NorthIn(nOut14_8), .SouthIn(nOut14_10), .EastIn(nOut15_9), .WestIn(nOut13_9), .ScanIn(nScanOut234), .ScanOut(nScanOut233), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_234 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_10), .NorthIn(nOut14_9), .SouthIn(nOut14_11), .EastIn(nOut15_10), .WestIn(nOut13_10), .ScanIn(nScanOut235), .ScanOut(nScanOut234), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_235 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_11), .NorthIn(nOut14_10), .SouthIn(nOut14_12), .EastIn(nOut15_11), .WestIn(nOut13_11), .ScanIn(nScanOut236), .ScanOut(nScanOut235), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_236 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_12), .NorthIn(nOut14_11), .SouthIn(nOut14_13), .EastIn(nOut15_12), .WestIn(nOut13_12), .ScanIn(nScanOut237), .ScanOut(nScanOut236), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_237 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_13), .NorthIn(nOut14_12), .SouthIn(nOut14_14), .EastIn(nOut15_13), .WestIn(nOut13_13), .ScanIn(nScanOut238), .ScanOut(nScanOut237), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_238 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut14_14), .NorthIn(nOut14_13), .SouthIn(nOut14_15), .EastIn(nOut15_14), .WestIn(nOut13_14), .ScanIn(nScanOut239), .ScanOut(nScanOut238), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_239 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut14_15), .ScanIn(nScanOut240), .ScanOut(nScanOut239), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_240 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_0), .ScanIn(nScanOut241), .ScanOut(nScanOut240), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_241 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_1), .ScanIn(nScanOut242), .ScanOut(nScanOut241), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_242 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_2), .ScanIn(nScanOut243), .ScanOut(nScanOut242), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_243 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_3), .ScanIn(nScanOut244), .ScanOut(nScanOut243), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_244 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_4), .ScanIn(nScanOut245), .ScanOut(nScanOut244), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_245 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_5), .ScanIn(nScanOut246), .ScanOut(nScanOut245), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_246 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_6), .ScanIn(nScanOut247), .ScanOut(nScanOut246), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_247 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_7), .ScanIn(nScanOut248), .ScanOut(nScanOut247), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_248 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_8), .ScanIn(nScanOut249), .ScanOut(nScanOut248), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_249 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_9), .ScanIn(nScanOut250), .ScanOut(nScanOut249), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_250 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_10), .ScanIn(nScanOut251), .ScanOut(nScanOut250), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_251 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_11), .ScanIn(nScanOut252), .ScanOut(nScanOut251), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_252 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_12), .ScanIn(nScanOut253), .ScanOut(nScanOut252), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_253 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_13), .ScanIn(nScanOut254), .ScanOut(nScanOut253), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_254 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_14), .ScanIn(nScanOut255), .ScanOut(nScanOut254), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_255 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut15_15), .ScanIn(nScanOut256), .ScanOut(nScanOut255), .ScanEnable(nScanEnable) );
Jacobi_Control #( 8, 7, 1, 1 ) U_Jacobi_Control ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Enable(nEnable), .ScanId(1'd0), .ScanEnable(nScanEnable), .ScanIn(nScanOut0), .ScanOut(nScanOut256) );

/*
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
