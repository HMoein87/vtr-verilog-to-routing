

/*
 *
 * RAW Benchmark Suite main defines
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */

`define GlobalDataWidth 32	    /* Global data bus width    */
`define GlobalAddrWidth 15	    /* Global address bus width */
				    /* Global data bus high impedance */
`define GlobalDataHighZ 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz 

/*
 * $Header: /projects/raw/cvsroot/benchmark/suites/jacobi/src/library.v,v 1.5 1997/08/09 05:57:41 jbabb Exp $
 *
 * Library for Jacobi benchmark
 *
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */



/*
 * This is the behavioral verilog library for this benchmark.
 * By convention, all module names start with the benchmark name.
 * All top-level modules must have the global connections:
 *   Clk, Reset, RD, WR, Addr, DataIn, DataOut
 * Modules may also have any number of local connections or
 * sub-modules without restriction.
 *
 */


/* The basic array node */

module Jacobi_Node (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		    ScanIn, ScanOut, ScanEnable,
		    Id, Enable, NorthIn, SouthIn, EastIn, WestIn, Out);
   
   parameter WIDTH    = 8,
	     IDWIDTH  = 8,
	     BOUNDARY = 0,
	     SCAN     = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   input			 ScanEnable;   


   /* local connections */
   
   input			 Enable;
   input [IDWIDTH-1:0]		 Id;
   input [WIDTH-1:0]		 NorthIn,SouthIn,EastIn,WestIn;
   output [WIDTH-1:0]		 Out;
   
   reg [WIDTH-1:0]		 Out;
   
   
   /* support reading of the node data value (non-scan only) */
   
   assign DataOut[`GlobalDataWidth-1:0] =
      (!SCAN && Addr[IDWIDTH-1:0] == Id) ? Out: `GlobalDataHighZ;


   /* support scan out of the node data value */

   assign ScanOut = SCAN ? Out: 0;

   
   always @(posedge Clk)
      begin	

	 
	 /* reset will initialize the entire array to zero */
	 
	 if (Reset)
	    Out=0;	 


	 /* support scan in */

	 else if (SCAN && ScanEnable)
	    Out=ScanIn[WIDTH-1:0];
	 

	 /* support writing of the node data value (non-scan only) */
	 
	 else if (!SCAN && WR && (Addr[IDWIDTH-1:0]==Id))
	    Out=DataIn[WIDTH-1:0];
	 

	 /* for non-boundary nodes, do the Jacobi computation when enabled */
	 
	 else if (!BOUNDARY && Enable)
	    Out=(NorthIn+SouthIn+EastIn+WestIn) >> 2;

      end
endmodule


/* 
 * A control module to count iterations.
 *
 * Writing to Address==ID will set a counter.
 *
 * The other Jacobi nodes will be enabled by this module when 
 * count is greater than zero.
 *
 * The counter will decrement every cycle down to zero.
 *
 * This module also handles scan control.
 */

module Jacobi_Control (Clk, Reset, RD, WR, Addr, DataIn, DataOut,
		       ScanIn, ScanOut, ScanEnable,
		       Id,ScanId,Enable);
   
   parameter WIDTH   = 8,
	     CWIDTH  = 8,
	     IDWIDTH = 8,
	     SCAN    = 1;
   
   
   /* global connections */
   
   input			 Clk,Reset,RD,WR;
   input [`GlobalAddrWidth-1:0]	 Addr;
   input [`GlobalDataWidth-1:0]	 DataIn;
   output [`GlobalDataWidth-1:0] DataOut;


   /* global connections for scan path (scan = 1) */

   input [IDWIDTH-1:0]		 ScanId;
   input [WIDTH-1:0]		 ScanIn;
   output [WIDTH-1:0]		 ScanOut;
   output			 ScanEnable;   


   /* local connections */
   
   input [IDWIDTH-1:0]		 Id;
   output			 Enable;
   
   
   /* a register for the counter and scan */

   reg [CWIDTH-1:0]		 count;
   reg [WIDTH-1:0]		 ScanReg;

   
   /* support writing scan input */

   assign ScanEnable=(SCAN && (RD || WR) && Addr[IDWIDTH-1:0]==ScanId);
   assign ScanOut= WR ? DataIn[WIDTH-1:0]: 0;


   /* support reading of the counter and scan output */

   assign DataOut[`GlobalDataWidth-1:0] =
      (Addr[IDWIDTH-1:0] == Id) ? count:
      (ScanEnable && RD) ? ScanReg: `GlobalDataHighZ;
   
   
   /* enable when count is active */
   
   assign Enable = !(count==0);

   
   always @(posedge Clk)
      begin

	 
	 /* store current scan output */

	 ScanReg=ScanIn;


	 /* Logic to reset, write, and decrement the counter */
	 
	 if (Reset)
	    count=0;
	 else if (WR && (Addr[IDWIDTH-1:0]==Id))
	    count=DataIn[CWIDTH-1:0];
	 else if(count) 
	    count=count-1;
      end
endmodule

/*
 *
 * RAW Benchmark Suite main module header
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


module main (
             Clk,
             Reset,
             RD,
             WR,
             Addr,
             DataIn,
             DataOut
            );

/* global connections */
input  Clk,Reset,RD,WR;
input  [`GlobalAddrWidth-1:0] Addr;
input  [`GlobalDataWidth-1:0] DataIn;
output [`GlobalDataWidth-1:0] DataOut;

wire [7:0] nOut0_0;
wire [7:0] nScanOut0;
wire [7:0] nOut0_1;
wire [7:0] nScanOut1;
wire [7:0] nOut0_2;
wire [7:0] nScanOut2;
wire [7:0] nOut0_3;
wire [7:0] nScanOut3;
wire [7:0] nOut0_4;
wire [7:0] nScanOut4;
wire [7:0] nOut0_5;
wire [7:0] nScanOut5;
wire [7:0] nOut0_6;
wire [7:0] nScanOut6;
wire [7:0] nOut0_7;
wire [7:0] nScanOut7;
wire [7:0] nOut1_0;
wire [7:0] nScanOut8;
wire [7:0] nOut1_1;
wire [7:0] nScanOut9;
wire [7:0] nOut1_2;
wire [7:0] nScanOut10;
wire [7:0] nOut1_3;
wire [7:0] nScanOut11;
wire [7:0] nOut1_4;
wire [7:0] nScanOut12;
wire [7:0] nOut1_5;
wire [7:0] nScanOut13;
wire [7:0] nOut1_6;
wire [7:0] nScanOut14;
wire [7:0] nOut1_7;
wire [7:0] nScanOut15;
wire [7:0] nOut2_0;
wire [7:0] nScanOut16;
wire [7:0] nOut2_1;
wire [7:0] nScanOut17;
wire [7:0] nOut2_2;
wire [7:0] nScanOut18;
wire [7:0] nOut2_3;
wire [7:0] nScanOut19;
wire [7:0] nOut2_4;
wire [7:0] nScanOut20;
wire [7:0] nOut2_5;
wire [7:0] nScanOut21;
wire [7:0] nOut2_6;
wire [7:0] nScanOut22;
wire [7:0] nOut2_7;
wire [7:0] nScanOut23;
wire [7:0] nOut3_0;
wire [7:0] nScanOut24;
wire [7:0] nOut3_1;
wire [7:0] nScanOut25;
wire [7:0] nOut3_2;
wire [7:0] nScanOut26;
wire [7:0] nOut3_3;
wire [7:0] nScanOut27;
wire [7:0] nOut3_4;
wire [7:0] nScanOut28;
wire [7:0] nOut3_5;
wire [7:0] nScanOut29;
wire [7:0] nOut3_6;
wire [7:0] nScanOut30;
wire [7:0] nOut3_7;
wire [7:0] nScanOut31;
wire [7:0] nOut4_0;
wire [7:0] nScanOut32;
wire [7:0] nOut4_1;
wire [7:0] nScanOut33;
wire [7:0] nOut4_2;
wire [7:0] nScanOut34;
wire [7:0] nOut4_3;
wire [7:0] nScanOut35;
wire [7:0] nOut4_4;
wire [7:0] nScanOut36;
wire [7:0] nOut4_5;
wire [7:0] nScanOut37;
wire [7:0] nOut4_6;
wire [7:0] nScanOut38;
wire [7:0] nOut4_7;
wire [7:0] nScanOut39;
wire [7:0] nOut5_0;
wire [7:0] nScanOut40;
wire [7:0] nOut5_1;
wire [7:0] nScanOut41;
wire [7:0] nOut5_2;
wire [7:0] nScanOut42;
wire [7:0] nOut5_3;
wire [7:0] nScanOut43;
wire [7:0] nOut5_4;
wire [7:0] nScanOut44;
wire [7:0] nOut5_5;
wire [7:0] nScanOut45;
wire [7:0] nOut5_6;
wire [7:0] nScanOut46;
wire [7:0] nOut5_7;
wire [7:0] nScanOut47;
wire [7:0] nOut6_0;
wire [7:0] nScanOut48;
wire [7:0] nOut6_1;
wire [7:0] nScanOut49;
wire [7:0] nOut6_2;
wire [7:0] nScanOut50;
wire [7:0] nOut6_3;
wire [7:0] nScanOut51;
wire [7:0] nOut6_4;
wire [7:0] nScanOut52;
wire [7:0] nOut6_5;
wire [7:0] nScanOut53;
wire [7:0] nOut6_6;
wire [7:0] nScanOut54;
wire [7:0] nOut6_7;
wire [7:0] nScanOut55;
wire [7:0] nOut7_0;
wire [7:0] nScanOut56;
wire [7:0] nOut7_1;
wire [7:0] nScanOut57;
wire [7:0] nOut7_2;
wire [7:0] nScanOut58;
wire [7:0] nOut7_3;
wire [7:0] nScanOut59;
wire [7:0] nOut7_4;
wire [7:0] nScanOut60;
wire [7:0] nOut7_5;
wire [7:0] nScanOut61;
wire [7:0] nOut7_6;
wire [7:0] nScanOut62;
wire [7:0] nOut7_7;
wire [7:0] nScanOut63;
wire [0:0] nEnable;
wire [0:0] nScanEnable;
wire [7:0] nScanOut64;
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_0 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_0), .ScanIn(nScanOut1), .ScanOut(nScanOut0), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_1 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_1), .ScanIn(nScanOut2), .ScanOut(nScanOut1), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_2 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_2), .ScanIn(nScanOut3), .ScanOut(nScanOut2), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_3 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_3), .ScanIn(nScanOut4), .ScanOut(nScanOut3), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_4 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_4), .ScanIn(nScanOut5), .ScanOut(nScanOut4), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_5 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_5), .ScanIn(nScanOut6), .ScanOut(nScanOut5), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_6 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_6), .ScanIn(nScanOut7), .ScanOut(nScanOut6), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_7 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut0_7), .ScanIn(nScanOut8), .ScanOut(nScanOut7), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_8 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_0), .ScanIn(nScanOut9), .ScanOut(nScanOut8), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_9 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_1), .NorthIn(nOut1_0), .SouthIn(nOut1_2), .EastIn(nOut2_1), .WestIn(nOut0_1), .ScanIn(nScanOut10), .ScanOut(nScanOut9), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_10 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_2), .NorthIn(nOut1_1), .SouthIn(nOut1_3), .EastIn(nOut2_2), .WestIn(nOut0_2), .ScanIn(nScanOut11), .ScanOut(nScanOut10), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_11 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_3), .NorthIn(nOut1_2), .SouthIn(nOut1_4), .EastIn(nOut2_3), .WestIn(nOut0_3), .ScanIn(nScanOut12), .ScanOut(nScanOut11), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_12 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_4), .NorthIn(nOut1_3), .SouthIn(nOut1_5), .EastIn(nOut2_4), .WestIn(nOut0_4), .ScanIn(nScanOut13), .ScanOut(nScanOut12), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_13 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_5), .NorthIn(nOut1_4), .SouthIn(nOut1_6), .EastIn(nOut2_5), .WestIn(nOut0_5), .ScanIn(nScanOut14), .ScanOut(nScanOut13), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_14 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut1_6), .NorthIn(nOut1_5), .SouthIn(nOut1_7), .EastIn(nOut2_6), .WestIn(nOut0_6), .ScanIn(nScanOut15), .ScanOut(nScanOut14), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_15 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut1_7), .ScanIn(nScanOut16), .ScanOut(nScanOut15), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_16 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_0), .ScanIn(nScanOut17), .ScanOut(nScanOut16), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_17 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_1), .NorthIn(nOut2_0), .SouthIn(nOut2_2), .EastIn(nOut3_1), .WestIn(nOut1_1), .ScanIn(nScanOut18), .ScanOut(nScanOut17), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_18 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_2), .NorthIn(nOut2_1), .SouthIn(nOut2_3), .EastIn(nOut3_2), .WestIn(nOut1_2), .ScanIn(nScanOut19), .ScanOut(nScanOut18), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_19 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_3), .NorthIn(nOut2_2), .SouthIn(nOut2_4), .EastIn(nOut3_3), .WestIn(nOut1_3), .ScanIn(nScanOut20), .ScanOut(nScanOut19), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_20 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_4), .NorthIn(nOut2_3), .SouthIn(nOut2_5), .EastIn(nOut3_4), .WestIn(nOut1_4), .ScanIn(nScanOut21), .ScanOut(nScanOut20), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_21 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_5), .NorthIn(nOut2_4), .SouthIn(nOut2_6), .EastIn(nOut3_5), .WestIn(nOut1_5), .ScanIn(nScanOut22), .ScanOut(nScanOut21), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_22 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut2_6), .NorthIn(nOut2_5), .SouthIn(nOut2_7), .EastIn(nOut3_6), .WestIn(nOut1_6), .ScanIn(nScanOut23), .ScanOut(nScanOut22), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_23 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut2_7), .ScanIn(nScanOut24), .ScanOut(nScanOut23), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_24 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_0), .ScanIn(nScanOut25), .ScanOut(nScanOut24), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_25 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_1), .NorthIn(nOut3_0), .SouthIn(nOut3_2), .EastIn(nOut4_1), .WestIn(nOut2_1), .ScanIn(nScanOut26), .ScanOut(nScanOut25), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_26 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_2), .NorthIn(nOut3_1), .SouthIn(nOut3_3), .EastIn(nOut4_2), .WestIn(nOut2_2), .ScanIn(nScanOut27), .ScanOut(nScanOut26), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_27 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_3), .NorthIn(nOut3_2), .SouthIn(nOut3_4), .EastIn(nOut4_3), .WestIn(nOut2_3), .ScanIn(nScanOut28), .ScanOut(nScanOut27), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_28 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_4), .NorthIn(nOut3_3), .SouthIn(nOut3_5), .EastIn(nOut4_4), .WestIn(nOut2_4), .ScanIn(nScanOut29), .ScanOut(nScanOut28), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_29 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_5), .NorthIn(nOut3_4), .SouthIn(nOut3_6), .EastIn(nOut4_5), .WestIn(nOut2_5), .ScanIn(nScanOut30), .ScanOut(nScanOut29), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_30 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut3_6), .NorthIn(nOut3_5), .SouthIn(nOut3_7), .EastIn(nOut4_6), .WestIn(nOut2_6), .ScanIn(nScanOut31), .ScanOut(nScanOut30), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_31 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut3_7), .ScanIn(nScanOut32), .ScanOut(nScanOut31), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_32 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_0), .ScanIn(nScanOut33), .ScanOut(nScanOut32), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_33 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_1), .NorthIn(nOut4_0), .SouthIn(nOut4_2), .EastIn(nOut5_1), .WestIn(nOut3_1), .ScanIn(nScanOut34), .ScanOut(nScanOut33), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_34 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_2), .NorthIn(nOut4_1), .SouthIn(nOut4_3), .EastIn(nOut5_2), .WestIn(nOut3_2), .ScanIn(nScanOut35), .ScanOut(nScanOut34), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_35 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_3), .NorthIn(nOut4_2), .SouthIn(nOut4_4), .EastIn(nOut5_3), .WestIn(nOut3_3), .ScanIn(nScanOut36), .ScanOut(nScanOut35), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_36 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_4), .NorthIn(nOut4_3), .SouthIn(nOut4_5), .EastIn(nOut5_4), .WestIn(nOut3_4), .ScanIn(nScanOut37), .ScanOut(nScanOut36), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_37 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_5), .NorthIn(nOut4_4), .SouthIn(nOut4_6), .EastIn(nOut5_5), .WestIn(nOut3_5), .ScanIn(nScanOut38), .ScanOut(nScanOut37), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_38 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut4_6), .NorthIn(nOut4_5), .SouthIn(nOut4_7), .EastIn(nOut5_6), .WestIn(nOut3_6), .ScanIn(nScanOut39), .ScanOut(nScanOut38), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_39 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut4_7), .ScanIn(nScanOut40), .ScanOut(nScanOut39), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_40 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_0), .ScanIn(nScanOut41), .ScanOut(nScanOut40), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_41 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_1), .NorthIn(nOut5_0), .SouthIn(nOut5_2), .EastIn(nOut6_1), .WestIn(nOut4_1), .ScanIn(nScanOut42), .ScanOut(nScanOut41), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_42 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_2), .NorthIn(nOut5_1), .SouthIn(nOut5_3), .EastIn(nOut6_2), .WestIn(nOut4_2), .ScanIn(nScanOut43), .ScanOut(nScanOut42), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_43 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_3), .NorthIn(nOut5_2), .SouthIn(nOut5_4), .EastIn(nOut6_3), .WestIn(nOut4_3), .ScanIn(nScanOut44), .ScanOut(nScanOut43), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_44 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_4), .NorthIn(nOut5_3), .SouthIn(nOut5_5), .EastIn(nOut6_4), .WestIn(nOut4_4), .ScanIn(nScanOut45), .ScanOut(nScanOut44), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_45 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_5), .NorthIn(nOut5_4), .SouthIn(nOut5_6), .EastIn(nOut6_5), .WestIn(nOut4_5), .ScanIn(nScanOut46), .ScanOut(nScanOut45), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_46 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut5_6), .NorthIn(nOut5_5), .SouthIn(nOut5_7), .EastIn(nOut6_6), .WestIn(nOut4_6), .ScanIn(nScanOut47), .ScanOut(nScanOut46), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_47 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut5_7), .ScanIn(nScanOut48), .ScanOut(nScanOut47), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_48 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_0), .ScanIn(nScanOut49), .ScanOut(nScanOut48), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_49 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_1), .NorthIn(nOut6_0), .SouthIn(nOut6_2), .EastIn(nOut7_1), .WestIn(nOut5_1), .ScanIn(nScanOut50), .ScanOut(nScanOut49), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_50 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_2), .NorthIn(nOut6_1), .SouthIn(nOut6_3), .EastIn(nOut7_2), .WestIn(nOut5_2), .ScanIn(nScanOut51), .ScanOut(nScanOut50), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_51 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_3), .NorthIn(nOut6_2), .SouthIn(nOut6_4), .EastIn(nOut7_3), .WestIn(nOut5_3), .ScanIn(nScanOut52), .ScanOut(nScanOut51), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_52 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_4), .NorthIn(nOut6_3), .SouthIn(nOut6_5), .EastIn(nOut7_4), .WestIn(nOut5_4), .ScanIn(nScanOut53), .ScanOut(nScanOut52), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_53 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_5), .NorthIn(nOut6_4), .SouthIn(nOut6_6), .EastIn(nOut7_5), .WestIn(nOut5_5), .ScanIn(nScanOut54), .ScanOut(nScanOut53), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 0, 1 ) U_Jacobi_Node_54 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Enable(nEnable), .Out(nOut6_6), .NorthIn(nOut6_5), .SouthIn(nOut6_7), .EastIn(nOut7_6), .WestIn(nOut5_6), .ScanIn(nScanOut55), .ScanOut(nScanOut54), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_55 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut6_7), .ScanIn(nScanOut56), .ScanOut(nScanOut55), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_56 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_0), .ScanIn(nScanOut57), .ScanOut(nScanOut56), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_57 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_1), .ScanIn(nScanOut58), .ScanOut(nScanOut57), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_58 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_2), .ScanIn(nScanOut59), .ScanOut(nScanOut58), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_59 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_3), .ScanIn(nScanOut60), .ScanOut(nScanOut59), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_60 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_4), .ScanIn(nScanOut61), .ScanOut(nScanOut60), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_61 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_5), .ScanIn(nScanOut62), .ScanOut(nScanOut61), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_62 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_6), .ScanIn(nScanOut63), .ScanOut(nScanOut62), .ScanEnable(nScanEnable) );
Jacobi_Node #( 8, 1, 1, 1 ) U_Jacobi_Node_63 ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd0), .Out(nOut7_7), .ScanIn(nScanOut64), .ScanOut(nScanOut63), .ScanEnable(nScanEnable) );
Jacobi_Control #( 8, 7, 1, 1 ) U_Jacobi_Control ( .Clk(Clk), .Reset(Reset), .RD(RD), .WR(WR), .Addr(Addr), .DataIn(DataIn), .DataOut(DataOut), .Id(1'd1), .Enable(nEnable), .ScanId(1'd0), .ScanEnable(nScanEnable), .ScanIn(nScanOut0), .ScanOut(nScanOut64) );

/*
 *
 * RAW Benchmark Suite main module trailer
 * 
 * Authors: Jonathan Babb           (jbabb@lcs.mit.edu)
 *
 * Copyright @ 1997 MIT Laboratory for Computer Science, Cambridge, MA 02129
 */


endmodule
